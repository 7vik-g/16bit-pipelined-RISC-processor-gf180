// This is the unpowered netlist.
module multiply_komal (Clock,
    Enable,
    done,
    reset,
    K,
    Result,
    X,
    Z);
 input Clock;
 input Enable;
 output done;
 input reset;
 input [2:0] K;
 output [16:0] Result;
 input [7:0] X;
 input [1:0] Z;

 wire \A[0][0] ;
 wire \A[0][1] ;
 wire \A[0][2] ;
 wire \A[0][3] ;
 wire \A[0][4] ;
 wire \A[0][5] ;
 wire \A[0][6] ;
 wire \A[0][7] ;
 wire \A[1][0] ;
 wire \A[1][1] ;
 wire \A[1][2] ;
 wire \A[1][3] ;
 wire \A[1][4] ;
 wire \A[1][5] ;
 wire \A[1][6] ;
 wire \A[1][7] ;
 wire \A[2][0] ;
 wire \A[2][1] ;
 wire \A[2][2] ;
 wire \A[2][3] ;
 wire \A[2][4] ;
 wire \A[2][5] ;
 wire \A[2][6] ;
 wire \A[2][7] ;
 wire \A[3][0] ;
 wire \A[3][1] ;
 wire \A[3][2] ;
 wire \A[3][3] ;
 wire \A[3][4] ;
 wire \A[3][5] ;
 wire \A[3][6] ;
 wire \A[3][7] ;
 wire \B[0][0] ;
 wire \B[0][1] ;
 wire \B[0][2] ;
 wire \B[0][3] ;
 wire \B[0][4] ;
 wire \B[0][5] ;
 wire \B[0][6] ;
 wire \B[0][7] ;
 wire \B[1][0] ;
 wire \B[1][1] ;
 wire \B[1][2] ;
 wire \B[1][3] ;
 wire \B[1][4] ;
 wire \B[1][5] ;
 wire \B[1][6] ;
 wire \B[1][7] ;
 wire \B[2][0] ;
 wire \B[2][1] ;
 wire \B[2][2] ;
 wire \B[2][3] ;
 wire \B[2][4] ;
 wire \B[2][5] ;
 wire \B[2][6] ;
 wire \B[2][7] ;
 wire \B[3][0] ;
 wire \B[3][1] ;
 wire \B[3][2] ;
 wire \B[3][3] ;
 wire \B[3][4] ;
 wire \B[3][5] ;
 wire \B[3][6] ;
 wire \B[3][7] ;
 wire \C[0][0] ;
 wire \C[0][10] ;
 wire \C[0][11] ;
 wire \C[0][12] ;
 wire \C[0][13] ;
 wire \C[0][14] ;
 wire \C[0][15] ;
 wire \C[0][16] ;
 wire \C[0][1] ;
 wire \C[0][2] ;
 wire \C[0][3] ;
 wire \C[0][4] ;
 wire \C[0][5] ;
 wire \C[0][6] ;
 wire \C[0][7] ;
 wire \C[0][8] ;
 wire \C[0][9] ;
 wire \C[1][0] ;
 wire \C[1][10] ;
 wire \C[1][11] ;
 wire \C[1][12] ;
 wire \C[1][13] ;
 wire \C[1][14] ;
 wire \C[1][15] ;
 wire \C[1][16] ;
 wire \C[1][1] ;
 wire \C[1][2] ;
 wire \C[1][3] ;
 wire \C[1][4] ;
 wire \C[1][5] ;
 wire \C[1][6] ;
 wire \C[1][7] ;
 wire \C[1][8] ;
 wire \C[1][9] ;
 wire \C[2][0] ;
 wire \C[2][10] ;
 wire \C[2][11] ;
 wire \C[2][12] ;
 wire \C[2][13] ;
 wire \C[2][14] ;
 wire \C[2][15] ;
 wire \C[2][16] ;
 wire \C[2][1] ;
 wire \C[2][2] ;
 wire \C[2][3] ;
 wire \C[2][4] ;
 wire \C[2][5] ;
 wire \C[2][6] ;
 wire \C[2][7] ;
 wire \C[2][8] ;
 wire \C[2][9] ;
 wire \C[3][0] ;
 wire \C[3][10] ;
 wire \C[3][11] ;
 wire \C[3][12] ;
 wire \C[3][13] ;
 wire \C[3][14] ;
 wire \C[3][15] ;
 wire \C[3][16] ;
 wire \C[3][1] ;
 wire \C[3][2] ;
 wire \C[3][3] ;
 wire \C[3][4] ;
 wire \C[3][5] ;
 wire \C[3][6] ;
 wire \C[3][7] ;
 wire \C[3][8] ;
 wire \C[3][9] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire clknet_0_Clock;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire clknet_3_0_0_Clock;
 wire clknet_3_1_0_Clock;
 wire clknet_3_2_0_Clock;
 wire clknet_3_3_0_Clock;
 wire clknet_3_4_0_Clock;
 wire clknet_3_5_0_Clock;
 wire clknet_3_6_0_Clock;
 wire clknet_3_7_0_Clock;
 wire clknet_4_0_0_Clock;
 wire clknet_4_1_0_Clock;
 wire clknet_4_2_0_Clock;
 wire clknet_4_3_0_Clock;
 wire clknet_4_4_0_Clock;
 wire clknet_4_5_0_Clock;
 wire clknet_4_6_0_Clock;
 wire clknet_4_7_0_Clock;
 wire clknet_4_8_0_Clock;
 wire clknet_4_9_0_Clock;
 wire clknet_4_10_0_Clock;
 wire clknet_4_11_0_Clock;
 wire clknet_4_12_0_Clock;
 wire clknet_4_13_0_Clock;
 wire clknet_4_14_0_Clock;
 wire clknet_4_15_0_Clock;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;

 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4277_ (.I(net1),
    .Z(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4278_ (.I(net3),
    .Z(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4279_ (.I(_2244_),
    .Z(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4280_ (.I(net2),
    .Z(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4281_ (.I(_2265_),
    .Z(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4282_ (.I(net4),
    .Z(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4283_ (.A1(_2233_),
    .A2(_2254_),
    .A3(_2276_),
    .A4(_2287_),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4284_ (.A1(\B[3][2] ),
    .A2(_2298_),
    .Z(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4285_ (.I(net1),
    .Z(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4286_ (.I(_2319_),
    .Z(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4287_ (.A1(_2330_),
    .A2(net7),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4288_ (.I(_2254_),
    .Z(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4289_ (.I(net2),
    .Z(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4290_ (.I(_2362_),
    .Z(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4291_ (.I(net4),
    .Z(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4292_ (.I(_2383_),
    .Z(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4293_ (.A1(_2352_),
    .A2(_2373_),
    .A3(_2394_),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4294_ (.A1(_2341_),
    .A2(_2405_),
    .ZN(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4295_ (.A1(_2308_),
    .A2(_2416_),
    .ZN(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4296_ (.I(_2427_),
    .ZN(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4297_ (.I(_2438_),
    .Z(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4298_ (.I(_2449_),
    .Z(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4299_ (.I(net1),
    .ZN(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4300_ (.I(_2470_),
    .Z(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4301_ (.I(_2481_),
    .Z(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4302_ (.I(_2383_),
    .Z(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4303_ (.I(_2503_),
    .Z(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4304_ (.A1(_2254_),
    .A2(_2276_),
    .ZN(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4305_ (.I(_2524_),
    .Z(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4306_ (.A1(_2492_),
    .A2(_2513_),
    .A3(_2534_),
    .B(\A[3][3] ),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _4307_ (.I(_2383_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4308_ (.I(_2556_),
    .Z(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4309_ (.I(_2567_),
    .Z(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4310_ (.A1(_2319_),
    .A2(net8),
    .Z(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4311_ (.I(_2589_),
    .Z(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4312_ (.I(net3),
    .Z(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4313_ (.A1(_2610_),
    .A2(_2362_),
    .Z(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4314_ (.I(_2621_),
    .Z(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4315_ (.A1(_2578_),
    .A2(_2599_),
    .A3(_2631_),
    .ZN(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4316_ (.I(net15),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4317_ (.A1(_2319_),
    .A2(_2652_),
    .ZN(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4318_ (.I(_2663_),
    .Z(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4319_ (.A1(_2545_),
    .A2(_2642_),
    .B(_2674_),
    .ZN(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4320_ (.I(_2685_),
    .Z(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4321_ (.I(_2695_),
    .Z(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4322_ (.I(_2706_),
    .Z(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4323_ (.A1(_2460_),
    .A2(_2717_),
    .Z(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4324_ (.I(_2470_),
    .Z(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4325_ (.I(_2737_),
    .Z(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4326_ (.I(_2394_),
    .Z(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4327_ (.I(_2524_),
    .Z(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4328_ (.A1(_2745_),
    .A2(_2755_),
    .A3(_2764_),
    .B(\A[3][2] ),
    .ZN(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4329_ (.I(_2556_),
    .Z(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4330_ (.I(_2786_),
    .Z(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4331_ (.I(net1),
    .Z(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4332_ (.A1(_2805_),
    .A2(net7),
    .Z(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4333_ (.I(_2816_),
    .Z(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4334_ (.I(_2621_),
    .Z(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4335_ (.A1(_2794_),
    .A2(_2826_),
    .A3(_2836_),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4336_ (.I(_2663_),
    .Z(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4337_ (.I(_2856_),
    .Z(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4338_ (.A1(_2775_),
    .A2(_2845_),
    .B(_2867_),
    .ZN(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4339_ (.I(_2878_),
    .Z(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4340_ (.I(_2589_),
    .Z(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4341_ (.A1(_2610_),
    .A2(_2362_),
    .A3(_2287_),
    .Z(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4342_ (.I(_2908_),
    .Z(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4343_ (.I(_2298_),
    .Z(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4344_ (.A1(_2897_),
    .A2(_2919_),
    .B1(_2930_),
    .B2(\B[3][3] ),
    .ZN(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4345_ (.I(_2941_),
    .ZN(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4346_ (.I(_2952_),
    .Z(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4347_ (.A1(_2889_),
    .A2(_2963_),
    .ZN(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4348_ (.A1(_2805_),
    .A2(net9),
    .Z(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4349_ (.A1(_2982_),
    .A2(_2908_),
    .B1(_2298_),
    .B2(\B[3][4] ),
    .ZN(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4350_ (.I(_2993_),
    .Z(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4351_ (.I(_3004_),
    .ZN(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4352_ (.I(_3015_),
    .Z(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4353_ (.I(_2737_),
    .Z(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4354_ (.I(_2503_),
    .Z(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4355_ (.A1(_3037_),
    .A2(_3048_),
    .A3(_2534_),
    .B(\A[3][1] ),
    .ZN(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4356_ (.I(_2786_),
    .Z(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4357_ (.A1(_2805_),
    .A2(net6),
    .Z(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4358_ (.A1(_3067_),
    .A2(_3078_),
    .A3(_2631_),
    .ZN(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4359_ (.I(_2856_),
    .Z(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4360_ (.A1(_3056_),
    .A2(_3089_),
    .B(_3100_),
    .ZN(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4361_ (.I(_3111_),
    .Z(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4362_ (.I(_3122_),
    .Z(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4363_ (.A1(_3026_),
    .A2(_3133_),
    .ZN(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4364_ (.A1(_2971_),
    .A2(_3144_),
    .Z(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4365_ (.A1(_2971_),
    .A2(_3144_),
    .ZN(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4366_ (.A1(_2727_),
    .A2(_3152_),
    .B(_3163_),
    .ZN(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4367_ (.I(_2330_),
    .Z(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4368_ (.A1(_3185_),
    .A2(net6),
    .ZN(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4369_ (.A1(\B[3][1] ),
    .A2(_2930_),
    .ZN(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4370_ (.A1(_3196_),
    .A2(_2405_),
    .B(_3207_),
    .ZN(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4371_ (.I(_3218_),
    .Z(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4372_ (.I(_3229_),
    .Z(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4373_ (.A1(_2745_),
    .A2(_3048_),
    .A3(_2534_),
    .B(\A[3][5] ),
    .ZN(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4374_ (.A1(_2805_),
    .A2(net10),
    .Z(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4375_ (.I(_3260_),
    .Z(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4376_ (.A1(_3067_),
    .A2(_3271_),
    .A3(_2631_),
    .ZN(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4377_ (.A1(_3249_),
    .A2(_3282_),
    .B(_3100_),
    .ZN(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4378_ (.I(_3293_),
    .Z(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4379_ (.I(_3304_),
    .Z(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4380_ (.I(_3315_),
    .Z(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4381_ (.A1(_3240_),
    .A2(_3326_),
    .ZN(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4382_ (.A1(_3174_),
    .A2(_3337_),
    .Z(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4383_ (.I(_2319_),
    .Z(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4384_ (.I(net5),
    .ZN(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4385_ (.A1(_3358_),
    .A2(_3369_),
    .ZN(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4386_ (.I(_3380_),
    .Z(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4387_ (.I(_2233_),
    .Z(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4388_ (.I(_3402_),
    .Z(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4389_ (.I(_3413_),
    .Z(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4390_ (.I(_3423_),
    .Z(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4391_ (.I(_2276_),
    .Z(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4392_ (.I(_2503_),
    .Z(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4393_ (.I(_3456_),
    .Z(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4394_ (.A1(_3434_),
    .A2(_2352_),
    .A3(_3445_),
    .A4(_3467_),
    .Z(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4395_ (.A1(_3391_),
    .A2(_2405_),
    .B1(_3478_),
    .B2(\B[3][0] ),
    .ZN(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4396_ (.I(_3488_),
    .ZN(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4397_ (.I(_3499_),
    .Z(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4398_ (.I(_3510_),
    .Z(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4399_ (.I(_2470_),
    .Z(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4400_ (.I(_3531_),
    .Z(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _4401_ (.A1(_3542_),
    .A2(_2755_),
    .A3(_2764_),
    .B(\A[3][6] ),
    .ZN(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _4402_ (.A1(_2330_),
    .A2(net11),
    .Z(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4403_ (.I(_3562_),
    .Z(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4404_ (.A1(_2794_),
    .A2(_2836_),
    .A3(_3572_),
    .ZN(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4405_ (.I(_2674_),
    .Z(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _4406_ (.A1(_3551_),
    .A2(_3583_),
    .B(_3593_),
    .ZN(_3604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4407_ (.I(_3604_),
    .Z(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4408_ (.I(_3615_),
    .Z(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4409_ (.I(_3625_),
    .Z(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4410_ (.I(_3636_),
    .Z(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4411_ (.I(_3646_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4412_ (.A1(_3174_),
    .A2(_3337_),
    .Z(_3662_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4413_ (.A1(_0056_),
    .A2(_0030_),
    .A3(_3662_),
    .ZN(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4414_ (.A1(_3347_),
    .A2(_3672_),
    .Z(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4415_ (.A1(_2481_),
    .A2(net15),
    .ZN(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4416_ (.I(_3691_),
    .Z(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4417_ (.I(_3701_),
    .Z(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4418_ (.I(\A[2][3] ),
    .ZN(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _4419_ (.I(_2244_),
    .ZN(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4420_ (.A1(_2737_),
    .A2(_3727_),
    .A3(_2373_),
    .A4(_2503_),
    .ZN(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4421_ (.I(_3735_),
    .Z(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4422_ (.A1(_3185_),
    .A2(net8),
    .ZN(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4423_ (.I(_2244_),
    .Z(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_8 _4424_ (.I(_2265_),
    .ZN(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 _4425_ (.I(_3747_),
    .Z(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4426_ (.A1(_3746_),
    .A2(_3748_),
    .A3(_2567_),
    .ZN(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4427_ (.I(_3749_),
    .Z(_3750_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _4428_ (.A1(_3718_),
    .A2(_3744_),
    .B1(_3745_),
    .B2(_3750_),
    .ZN(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4429_ (.I(\B[1][2] ),
    .ZN(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4430_ (.A1(_2737_),
    .A2(_3746_),
    .A3(_3747_),
    .A4(_2567_),
    .ZN(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4431_ (.I(_3753_),
    .Z(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4432_ (.A1(_3727_),
    .A2(_2373_),
    .A3(_2394_),
    .ZN(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4433_ (.I(_3755_),
    .Z(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4434_ (.A1(_3752_),
    .A2(_3754_),
    .B1(_2341_),
    .B2(_3756_),
    .ZN(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4435_ (.A1(_3709_),
    .A2(_3751_),
    .A3(_3757_),
    .ZN(_3758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4436_ (.I(_3691_),
    .Z(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4437_ (.I(_3759_),
    .Z(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4438_ (.I(_3760_),
    .Z(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4439_ (.I(_3761_),
    .Z(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4440_ (.I(\B[1][1] ),
    .ZN(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4441_ (.I(_3753_),
    .Z(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4442_ (.I(_3755_),
    .Z(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _4443_ (.A1(_3763_),
    .A2(_3764_),
    .B1(_3196_),
    .B2(_3765_),
    .ZN(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4444_ (.I(_3766_),
    .Z(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4445_ (.I(\A[2][2] ),
    .ZN(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4446_ (.I(_3735_),
    .Z(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4447_ (.I(_3749_),
    .Z(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4448_ (.A1(_3768_),
    .A2(_3769_),
    .B1(_2341_),
    .B2(_3770_),
    .ZN(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4449_ (.I(_3771_),
    .Z(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4450_ (.I(_3772_),
    .Z(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4451_ (.A1(_3762_),
    .A2(_3767_),
    .A3(_3773_),
    .ZN(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4452_ (.I(_2856_),
    .Z(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4453_ (.I(_3775_),
    .Z(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4454_ (.I(_3776_),
    .Z(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4455_ (.I(_3777_),
    .Z(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4456_ (.I(_3727_),
    .Z(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4457_ (.A1(_3402_),
    .A2(_3779_),
    .A3(_3445_),
    .A4(_2513_),
    .ZN(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4458_ (.I(_3780_),
    .Z(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4459_ (.I(_2556_),
    .Z(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4460_ (.A1(_2352_),
    .A2(_3748_),
    .A3(_3782_),
    .ZN(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4461_ (.I(_3783_),
    .Z(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4462_ (.A1(\B[1][2] ),
    .A2(_3781_),
    .B1(_2826_),
    .B2(_3784_),
    .ZN(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4463_ (.I(_3785_),
    .Z(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4464_ (.A1(_3402_),
    .A2(_2352_),
    .A3(_3748_),
    .A4(_3782_),
    .ZN(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4465_ (.A1(_3779_),
    .A2(_3445_),
    .A3(_2513_),
    .ZN(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4466_ (.A1(\A[2][2] ),
    .A2(_3787_),
    .B1(_2826_),
    .B2(_3788_),
    .ZN(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4467_ (.I(_3789_),
    .Z(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4468_ (.A1(_3778_),
    .A2(_3786_),
    .A3(_3790_),
    .ZN(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4469_ (.I(_3775_),
    .Z(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4470_ (.I(_3792_),
    .Z(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4471_ (.I(_3793_),
    .Z(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4472_ (.A1(\A[2][3] ),
    .A2(_3787_),
    .B1(_2897_),
    .B2(_3788_),
    .ZN(_3795_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4473_ (.I(_3795_),
    .Z(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4474_ (.I(_3078_),
    .Z(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4475_ (.A1(\B[1][1] ),
    .A2(_3781_),
    .B1(_3797_),
    .B2(_3784_),
    .ZN(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4476_ (.I(_3798_),
    .Z(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4477_ (.A1(_3794_),
    .A2(_3796_),
    .A3(_3799_),
    .ZN(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4478_ (.A1(_3758_),
    .A2(_3774_),
    .B1(_3791_),
    .B2(_3800_),
    .ZN(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4479_ (.A1(_2233_),
    .A2(net9),
    .ZN(_3802_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4480_ (.I(\A[2][4] ),
    .ZN(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4481_ (.A1(_3802_),
    .A2(_3750_),
    .B1(_3744_),
    .B2(_3803_),
    .ZN(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4482_ (.I(_3804_),
    .Z(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4483_ (.I(_3805_),
    .Z(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _4484_ (.A1(\B[1][0] ),
    .A2(_3754_),
    .B1(_3380_),
    .B2(_3756_),
    .C(_3701_),
    .ZN(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4485_ (.I(_3807_),
    .ZN(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4486_ (.I(_3808_),
    .Z(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4487_ (.A1(_3806_),
    .A2(_3809_),
    .ZN(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4488_ (.A1(_3758_),
    .A2(_3774_),
    .B1(_3801_),
    .B2(_3810_),
    .ZN(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _4489_ (.A1(\A[2][0] ),
    .A2(_3744_),
    .B1(_3391_),
    .B2(_3750_),
    .C(_3701_),
    .ZN(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _4490_ (.I(_3812_),
    .ZN(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4491_ (.I(_3813_),
    .Z(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4492_ (.I(\B[1][3] ),
    .ZN(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4493_ (.A1(_3815_),
    .A2(_3754_),
    .B1(_3745_),
    .B2(_3756_),
    .ZN(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4494_ (.I(_3816_),
    .Z(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4495_ (.I(_3817_),
    .Z(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4496_ (.I(_2982_),
    .Z(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4497_ (.A1(\B[1][4] ),
    .A2(_3781_),
    .B1(_3819_),
    .B2(_3784_),
    .ZN(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4498_ (.I(_2867_),
    .Z(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4499_ (.I(_3821_),
    .Z(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4500_ (.A1(\A[2][1] ),
    .A2(_3787_),
    .B1(_3797_),
    .B2(_3788_),
    .ZN(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4501_ (.I(_3823_),
    .Z(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4502_ (.A1(_3820_),
    .A2(_3822_),
    .A3(_3824_),
    .ZN(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4503_ (.A1(_3814_),
    .A2(_3818_),
    .A3(_3825_),
    .ZN(_3826_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4504_ (.A1(_3709_),
    .A2(_3766_),
    .A3(_3804_),
    .ZN(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4505_ (.I(\A[2][5] ),
    .ZN(_3828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4506_ (.A1(_3185_),
    .A2(net10),
    .ZN(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4507_ (.A1(_3828_),
    .A2(_3769_),
    .B1(_3829_),
    .B2(_3770_),
    .ZN(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4508_ (.I(_3830_),
    .Z(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4509_ (.I(_3808_),
    .Z(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4510_ (.A1(_3831_),
    .A2(_3832_),
    .ZN(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4511_ (.A1(_3758_),
    .A2(_3827_),
    .A3(_3833_),
    .Z(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4512_ (.A1(_3826_),
    .A2(_3834_),
    .Z(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4513_ (.A1(_3826_),
    .A2(_3834_),
    .ZN(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4514_ (.A1(_3811_),
    .A2(_3835_),
    .B(_3836_),
    .ZN(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4515_ (.A1(_3037_),
    .A2(_3048_),
    .A3(_2534_),
    .B(\A[3][4] ),
    .ZN(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4516_ (.A1(_3067_),
    .A2(_2982_),
    .A3(_2631_),
    .ZN(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4517_ (.A1(_3838_),
    .A2(_3839_),
    .B(_3775_),
    .ZN(_3840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4518_ (.I(_3840_),
    .Z(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4519_ (.I(_3841_),
    .Z(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4520_ (.A1(_2449_),
    .A2(_3842_),
    .Z(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4521_ (.I(_3015_),
    .Z(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4522_ (.I(_2695_),
    .Z(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4523_ (.A1(_3844_),
    .A2(_3845_),
    .ZN(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4524_ (.A1(_2971_),
    .A2(_3846_),
    .ZN(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4525_ (.I(_2889_),
    .Z(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4526_ (.I(_2963_),
    .Z(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4527_ (.A1(_3848_),
    .A2(_3026_),
    .B1(_2706_),
    .B2(_3849_),
    .ZN(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4528_ (.A1(_3847_),
    .A2(_3850_),
    .ZN(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4529_ (.A1(_3843_),
    .A2(_3851_),
    .ZN(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4530_ (.I(_2481_),
    .Z(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4531_ (.I(_3853_),
    .Z(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4532_ (.I(\A[3][0] ),
    .ZN(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4533_ (.A1(_3854_),
    .A2(_3467_),
    .A3(_2764_),
    .B(_3855_),
    .ZN(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4534_ (.A1(_3413_),
    .A2(_2794_),
    .A3(_3369_),
    .A4(_2836_),
    .ZN(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4535_ (.A1(_3760_),
    .A2(_3856_),
    .A3(_3857_),
    .ZN(_3858_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4536_ (.I(_3858_),
    .ZN(_3859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4537_ (.I(_3859_),
    .Z(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _4538_ (.A1(_3260_),
    .A2(_2919_),
    .B1(_2298_),
    .B2(\B[3][5] ),
    .ZN(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4539_ (.I(_3861_),
    .ZN(_3862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4540_ (.I(_3862_),
    .Z(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4541_ (.I(_3863_),
    .Z(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4542_ (.A1(_3860_),
    .A2(_3864_),
    .ZN(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4543_ (.A1(\B[3][6] ),
    .A2(_2930_),
    .B1(_3562_),
    .B2(_2919_),
    .ZN(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4544_ (.I(_3866_),
    .ZN(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4545_ (.A1(_3867_),
    .A2(_3122_),
    .ZN(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4546_ (.A1(_3865_),
    .A2(_3868_),
    .ZN(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4547_ (.I(_3860_),
    .Z(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4548_ (.I(_3870_),
    .Z(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4549_ (.I(_3867_),
    .Z(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4550_ (.I(_3872_),
    .Z(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4551_ (.I(_3873_),
    .Z(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4552_ (.I(_3122_),
    .Z(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4553_ (.I(_3875_),
    .Z(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4554_ (.I(_3864_),
    .Z(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4555_ (.A1(_3871_),
    .A2(_3874_),
    .B1(_3876_),
    .B2(_3877_),
    .ZN(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4556_ (.A1(_3869_),
    .A2(_3878_),
    .Z(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4557_ (.A1(_3852_),
    .A2(_3879_),
    .ZN(_3880_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4558_ (.A1(_3852_),
    .A2(_3879_),
    .Z(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4559_ (.I(_3870_),
    .Z(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4560_ (.I(_3877_),
    .Z(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4561_ (.I(_3883_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4562_ (.A1(_2727_),
    .A2(_3152_),
    .Z(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4563_ (.A1(_3882_),
    .A2(_0061_),
    .A3(_3884_),
    .ZN(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4564_ (.A1(_3837_),
    .A2(_3852_),
    .A3(_3879_),
    .Z(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4565_ (.A1(_3837_),
    .A2(_3880_),
    .A3(_3881_),
    .B1(_3885_),
    .B2(_3886_),
    .ZN(_3887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4566_ (.I(_3499_),
    .Z(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4567_ (.I(_3888_),
    .Z(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4568_ (.I(_2745_),
    .Z(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4569_ (.A1(_3890_),
    .A2(_3467_),
    .A3(_2764_),
    .B(\A[3][7] ),
    .ZN(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4570_ (.I(_3067_),
    .Z(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4571_ (.A1(_3358_),
    .A2(net12),
    .Z(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4572_ (.I(_3893_),
    .Z(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4573_ (.A1(_3892_),
    .A2(_2836_),
    .A3(_3894_),
    .ZN(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4574_ (.A1(_3891_),
    .A2(_3895_),
    .B(_3821_),
    .ZN(_3896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4575_ (.I(_3896_),
    .Z(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4576_ (.I(_3897_),
    .Z(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4577_ (.I(_3898_),
    .Z(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4578_ (.I(_3899_),
    .Z(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4579_ (.A1(_3889_),
    .A2(_3900_),
    .ZN(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4580_ (.A1(_3843_),
    .A2(_3851_),
    .B(_3847_),
    .ZN(_3902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4581_ (.I(_3229_),
    .Z(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4582_ (.I(_3903_),
    .Z(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4583_ (.I(_3636_),
    .Z(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4584_ (.A1(_3904_),
    .A2(_3905_),
    .ZN(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4585_ (.A1(_3902_),
    .A2(_3906_),
    .Z(_3907_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4586_ (.A1(_3901_),
    .A2(_3907_),
    .ZN(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4587_ (.A1(_3887_),
    .A2(_3908_),
    .ZN(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4588_ (.A1(_3887_),
    .A2(_3908_),
    .ZN(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4589_ (.A1(_3682_),
    .A2(_3909_),
    .B(_3910_),
    .ZN(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4590_ (.A1(_3682_),
    .A2(_3909_),
    .Z(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4591_ (.A1(_3885_),
    .A2(_3886_),
    .ZN(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4592_ (.A1(_3811_),
    .A2(_3835_),
    .ZN(_3914_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4593_ (.I(\B[1][4] ),
    .ZN(_3915_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4594_ (.A1(_3915_),
    .A2(_3753_),
    .B1(_3802_),
    .B2(_3755_),
    .ZN(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4595_ (.I(_3916_),
    .Z(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4596_ (.A1(_3917_),
    .A2(_3814_),
    .ZN(_3918_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4597_ (.I(\A[2][1] ),
    .ZN(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4598_ (.A1(_3919_),
    .A2(_3744_),
    .B1(_3196_),
    .B2(_3750_),
    .ZN(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4599_ (.I(_3920_),
    .Z(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4600_ (.I(_3921_),
    .Z(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4601_ (.A1(_3762_),
    .A2(_3922_),
    .A3(_3817_),
    .ZN(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4602_ (.A1(_3918_),
    .A2(_3923_),
    .ZN(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4603_ (.I(net15),
    .Z(_3925_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4604_ (.I(_3925_),
    .Z(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4605_ (.A1(_3423_),
    .A2(_3926_),
    .ZN(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4606_ (.I(_3927_),
    .Z(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4607_ (.I(_3928_),
    .Z(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4608_ (.A1(\C[3][4] ),
    .A2(_3826_),
    .A3(_3924_),
    .A4(_3929_),
    .Z(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4609_ (.I(_3916_),
    .Z(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4610_ (.A1(_3931_),
    .A2(_3761_),
    .A3(_3921_),
    .ZN(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4611_ (.I(\B[1][5] ),
    .ZN(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4612_ (.A1(_3933_),
    .A2(_3754_),
    .B1(_3829_),
    .B2(_3756_),
    .ZN(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4613_ (.A1(_3813_),
    .A2(_3934_),
    .ZN(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4614_ (.A1(\B[1][3] ),
    .A2(_3781_),
    .B1(_2897_),
    .B2(_3784_),
    .ZN(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4615_ (.I(_3789_),
    .Z(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4616_ (.A1(_3822_),
    .A2(_3936_),
    .A3(_3937_),
    .ZN(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4617_ (.A1(_3932_),
    .A2(_3935_),
    .A3(_3938_),
    .Z(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4618_ (.A1(\C[3][5] ),
    .A2(_3928_),
    .ZN(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4619_ (.A1(_3939_),
    .A2(_3940_),
    .ZN(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4620_ (.A1(_3930_),
    .A2(_3941_),
    .ZN(_3942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4621_ (.A1(_3930_),
    .A2(_3941_),
    .ZN(_3943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4622_ (.A1(_3914_),
    .A2(_3942_),
    .B(_3943_),
    .ZN(_3944_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4623_ (.A1(\C[3][5] ),
    .A2(_3929_),
    .A3(_3939_),
    .ZN(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4624_ (.I(_2856_),
    .Z(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4625_ (.I(_3946_),
    .Z(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4626_ (.I(_3947_),
    .Z(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4627_ (.A1(\B[1][5] ),
    .A2(_3780_),
    .B1(_3271_),
    .B2(_3783_),
    .ZN(_3949_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4628_ (.I(_3949_),
    .Z(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4629_ (.A1(_3948_),
    .A2(_3937_),
    .A3(_3950_),
    .ZN(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4630_ (.I(_3761_),
    .Z(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4631_ (.I(_3771_),
    .Z(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4632_ (.A1(_3931_),
    .A2(_3952_),
    .A3(_3953_),
    .ZN(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4633_ (.I(_3709_),
    .Z(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4634_ (.I(_3920_),
    .Z(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4635_ (.I(_3934_),
    .Z(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4636_ (.A1(_3955_),
    .A2(_3956_),
    .A3(_3957_),
    .ZN(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4637_ (.A1(_3825_),
    .A2(_3951_),
    .B1(_3954_),
    .B2(_3958_),
    .ZN(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4638_ (.I(_3946_),
    .Z(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4639_ (.I(_3960_),
    .Z(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4640_ (.I(_3936_),
    .Z(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4641_ (.A1(_3961_),
    .A2(_3962_),
    .A3(_3796_),
    .ZN(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4642_ (.I(_3813_),
    .Z(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4643_ (.I(_3964_),
    .Z(_3965_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4644_ (.I(\B[1][6] ),
    .ZN(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4645_ (.A1(_3413_),
    .A2(net11),
    .ZN(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4646_ (.A1(_3966_),
    .A2(_3764_),
    .B1(_3967_),
    .B2(_3765_),
    .ZN(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4647_ (.I(_3968_),
    .Z(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4648_ (.A1(_3965_),
    .A2(_3969_),
    .ZN(_3970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4649_ (.I(_3854_),
    .Z(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4650_ (.I(_3971_),
    .Z(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4651_ (.I(_3972_),
    .Z(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4652_ (.I(_2652_),
    .Z(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4653_ (.I(_3974_),
    .Z(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4654_ (.I(_3975_),
    .Z(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4655_ (.A1(_3973_),
    .A2(_3976_),
    .A3(\C[3][6] ),
    .ZN(_3977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4656_ (.I(_3812_),
    .Z(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4657_ (.I(_3978_),
    .Z(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4658_ (.A1(\B[1][6] ),
    .A2(_3780_),
    .B1(_3572_),
    .B2(_3783_),
    .ZN(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4659_ (.I(_3980_),
    .Z(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4660_ (.I(_3890_),
    .Z(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4661_ (.I(_3982_),
    .Z(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4662_ (.A1(_3983_),
    .A2(\C[3][6] ),
    .ZN(_3984_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4663_ (.A1(_3979_),
    .A2(_3981_),
    .A3(_3984_),
    .ZN(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4664_ (.A1(_3970_),
    .A2(_3977_),
    .B(_3985_),
    .ZN(_3986_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4665_ (.A1(_3959_),
    .A2(_3963_),
    .A3(_3986_),
    .ZN(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4666_ (.A1(_3945_),
    .A2(_3987_),
    .Z(_3988_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4667_ (.A1(_3758_),
    .A2(_3827_),
    .Z(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4668_ (.I(_2663_),
    .Z(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4669_ (.I(_3990_),
    .Z(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4670_ (.I(_3991_),
    .Z(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4671_ (.I(_3992_),
    .Z(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4672_ (.A1(_3993_),
    .A2(_3786_),
    .ZN(_3994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4673_ (.I(_3994_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4674_ (.A1(_3800_),
    .A2(_0042_),
    .A3(_3806_),
    .ZN(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4675_ (.A1(_3989_),
    .A2(_3833_),
    .B(_3995_),
    .ZN(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4676_ (.I(_3964_),
    .Z(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4677_ (.I(_3934_),
    .Z(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4678_ (.I(_3998_),
    .Z(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4679_ (.A1(_3997_),
    .A2(_3825_),
    .A3(_3999_),
    .ZN(_4000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4680_ (.I(_3820_),
    .Z(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4681_ (.I(_3823_),
    .Z(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4682_ (.I(_3949_),
    .Z(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4683_ (.A1(_4001_),
    .A2(_3778_),
    .A3(_4002_),
    .B1(_4003_),
    .B2(_3979_),
    .ZN(_4004_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4684_ (.A1(_3918_),
    .A2(_3958_),
    .B(_4004_),
    .C(_3938_),
    .ZN(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4685_ (.A1(_4000_),
    .A2(_4005_),
    .ZN(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4686_ (.I(_3757_),
    .Z(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4687_ (.A1(_3952_),
    .A2(_4007_),
    .A3(_3805_),
    .ZN(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4688_ (.I(_3766_),
    .Z(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4689_ (.I(_3830_),
    .Z(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4690_ (.A1(_3952_),
    .A2(_4009_),
    .A3(_4010_),
    .ZN(_4011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4691_ (.I(_3832_),
    .Z(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4692_ (.I(\A[2][6] ),
    .ZN(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4693_ (.A1(_4013_),
    .A2(_3769_),
    .B1(_3967_),
    .B2(_3770_),
    .ZN(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4694_ (.I(_4014_),
    .Z(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4695_ (.A1(_4012_),
    .A2(_4015_),
    .ZN(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4696_ (.A1(_4008_),
    .A2(_4011_),
    .A3(_4016_),
    .Z(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4697_ (.A1(_3996_),
    .A2(_4006_),
    .A3(_4017_),
    .ZN(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4698_ (.A1(_3988_),
    .A2(_4018_),
    .Z(_4019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4699_ (.A1(_3944_),
    .A2(_4019_),
    .ZN(_4020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4700_ (.A1(_3944_),
    .A2(_4019_),
    .ZN(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4701_ (.A1(_3913_),
    .A2(_4020_),
    .B(_4021_),
    .ZN(_4022_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4702_ (.A1(_4000_),
    .A2(_4005_),
    .A3(_4017_),
    .ZN(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4703_ (.A1(_4000_),
    .A2(_4005_),
    .B(_4017_),
    .ZN(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4704_ (.A1(_3996_),
    .A2(_4023_),
    .B(_4024_),
    .ZN(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4705_ (.I(_3304_),
    .Z(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4706_ (.A1(_2449_),
    .A2(_4026_),
    .ZN(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4707_ (.A1(_3841_),
    .A2(_3849_),
    .ZN(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4708_ (.A1(_3846_),
    .A2(_4028_),
    .Z(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4709_ (.A1(_4027_),
    .A2(_4029_),
    .Z(_4030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4710_ (.I(_2878_),
    .Z(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4711_ (.A1(_4031_),
    .A2(_3863_),
    .ZN(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4712_ (.I(_3858_),
    .Z(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4713_ (.A1(\B[3][7] ),
    .A2(_2930_),
    .B1(_3893_),
    .B2(_2919_),
    .ZN(_4034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4714_ (.I(_4034_),
    .Z(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4715_ (.A1(_4033_),
    .A2(_4035_),
    .ZN(_4036_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4716_ (.A1(_3868_),
    .A2(_4032_),
    .A3(_4036_),
    .Z(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4717_ (.A1(_3869_),
    .A2(_4037_),
    .ZN(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4718_ (.A1(_4030_),
    .A2(_4038_),
    .ZN(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4719_ (.A1(_4025_),
    .A2(_4039_),
    .Z(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4720_ (.A1(_3880_),
    .A2(_4040_),
    .Z(_4041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4721_ (.A1(_3945_),
    .A2(_3987_),
    .ZN(_4042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4722_ (.A1(_3988_),
    .A2(_4018_),
    .B(_4042_),
    .ZN(_4043_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4723_ (.A1(_3952_),
    .A2(_3953_),
    .A3(_3957_),
    .ZN(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4724_ (.I(_3947_),
    .Z(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4725_ (.A1(_3820_),
    .A2(_4045_),
    .A3(_3937_),
    .ZN(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4726_ (.A1(_3993_),
    .A2(_4002_),
    .A3(_3950_),
    .ZN(_4047_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _4727_ (.A1(_3932_),
    .A2(_4044_),
    .B1(_4046_),
    .B2(_4047_),
    .C(_3963_),
    .ZN(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4728_ (.A1(_3959_),
    .A2(_3963_),
    .Z(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4729_ (.A1(_4048_),
    .A2(_4049_),
    .A3(_3986_),
    .ZN(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4730_ (.A1(_4008_),
    .A2(_4011_),
    .Z(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4731_ (.A1(_4008_),
    .A2(_4011_),
    .Z(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4732_ (.A1(_4051_),
    .A2(_4016_),
    .B(_4052_),
    .ZN(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4733_ (.A1(_3825_),
    .A2(_3951_),
    .ZN(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4734_ (.A1(_4054_),
    .A2(_4048_),
    .ZN(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4735_ (.I(_4014_),
    .Z(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4736_ (.A1(_3955_),
    .A2(_4009_),
    .A3(_4056_),
    .ZN(_4057_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4737_ (.A1(_3955_),
    .A2(_4007_),
    .A3(_3831_),
    .ZN(_4058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4738_ (.I(\A[2][7] ),
    .ZN(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4739_ (.A1(_3423_),
    .A2(net12),
    .ZN(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4740_ (.A1(_4059_),
    .A2(_3769_),
    .B1(_4060_),
    .B2(_3770_),
    .ZN(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4741_ (.I(_4061_),
    .Z(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4742_ (.A1(_4012_),
    .A2(_4062_),
    .ZN(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4743_ (.A1(_4057_),
    .A2(_4058_),
    .A3(_4063_),
    .Z(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4744_ (.A1(_4053_),
    .A2(_4055_),
    .A3(_4064_),
    .ZN(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4745_ (.I(_3821_),
    .Z(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4746_ (.I(_3795_),
    .Z(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4747_ (.A1(_4066_),
    .A2(_4067_),
    .A3(_3950_),
    .ZN(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4748_ (.I(_3917_),
    .Z(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4749_ (.I(_3955_),
    .Z(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4750_ (.I(_3751_),
    .Z(_4071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4751_ (.I(_4071_),
    .Z(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4752_ (.I(_4072_),
    .Z(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4753_ (.A1(_4069_),
    .A2(_4070_),
    .A3(_4073_),
    .ZN(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4754_ (.A1(_4046_),
    .A2(_4068_),
    .B1(_4074_),
    .B2(_4044_),
    .ZN(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4755_ (.I(_3818_),
    .Z(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4756_ (.I(_3788_),
    .Z(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4757_ (.I(_3787_),
    .Z(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4758_ (.A1(_3819_),
    .A2(_4077_),
    .B1(_4078_),
    .B2(\A[2][4] ),
    .ZN(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4759_ (.I(_4079_),
    .Z(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4760_ (.A1(_3778_),
    .A2(_4080_),
    .ZN(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4761_ (.I(_4081_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4762_ (.A1(_4076_),
    .A2(_0020_),
    .ZN(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4763_ (.A1(_4075_),
    .A2(_4082_),
    .Z(_4083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4764_ (.I(\B[1][7] ),
    .ZN(_4084_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4765_ (.A1(_4084_),
    .A2(_3764_),
    .B1(_4060_),
    .B2(_3765_),
    .ZN(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4766_ (.A1(_3983_),
    .A2(\C[3][7] ),
    .A3(_3964_),
    .A4(_4085_),
    .ZN(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4767_ (.I(_3925_),
    .Z(_4087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4768_ (.I(_4087_),
    .Z(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4769_ (.I(_3542_),
    .Z(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4770_ (.I(_4089_),
    .Z(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4771_ (.A1(_4090_),
    .A2(\C[3][7] ),
    .ZN(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4772_ (.A1(\B[1][7] ),
    .A2(_3780_),
    .B1(_3893_),
    .B2(_3783_),
    .ZN(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4773_ (.I(_4092_),
    .Z(_4093_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4774_ (.A1(_4088_),
    .A2(_4091_),
    .B1(_4093_),
    .B2(_3978_),
    .ZN(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4775_ (.A1(_4086_),
    .A2(_4094_),
    .Z(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4776_ (.I(_3980_),
    .Z(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4777_ (.A1(_3961_),
    .A2(_3824_),
    .A3(_4096_),
    .ZN(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4778_ (.A1(_3985_),
    .A2(_4095_),
    .A3(_4097_),
    .ZN(_4098_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4779_ (.A1(_4083_),
    .A2(_4098_),
    .ZN(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4780_ (.A1(_4050_),
    .A2(_4065_),
    .A3(_4099_),
    .ZN(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4781_ (.A1(_4043_),
    .A2(_4100_),
    .Z(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4782_ (.A1(_4041_),
    .A2(_4101_),
    .Z(_4102_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4783_ (.A1(_4022_),
    .A2(_4102_),
    .Z(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4784_ (.A1(_4022_),
    .A2(_4102_),
    .Z(_4104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4785_ (.A1(_3912_),
    .A2(_4103_),
    .B(_4104_),
    .ZN(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4786_ (.A1(_3902_),
    .A2(_3906_),
    .Z(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4787_ (.I(_3899_),
    .Z(_4107_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4788_ (.A1(_0056_),
    .A2(_4107_),
    .A3(_3907_),
    .ZN(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4789_ (.A1(_4106_),
    .A2(_4108_),
    .Z(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4790_ (.A1(_4025_),
    .A2(_4039_),
    .ZN(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4791_ (.A1(_3880_),
    .A2(_4040_),
    .B(_4110_),
    .ZN(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4792_ (.I(_2438_),
    .Z(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4793_ (.I(_4112_),
    .Z(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4794_ (.I(_4113_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4795_ (.I(_3326_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4796_ (.A1(_0058_),
    .A2(_0029_),
    .A3(_4029_),
    .ZN(_4114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4797_ (.A1(_3846_),
    .A2(_4028_),
    .B(_4114_),
    .ZN(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4798_ (.I(_3903_),
    .Z(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4799_ (.I(_4116_),
    .Z(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4800_ (.A1(_4107_),
    .A2(_4117_),
    .ZN(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4801_ (.A1(_4111_),
    .A2(_4115_),
    .A3(_4118_),
    .ZN(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4802_ (.A1(_4109_),
    .A2(_4119_),
    .Z(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4803_ (.A1(_4043_),
    .A2(_4100_),
    .ZN(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4804_ (.A1(_4041_),
    .A2(_4101_),
    .B(_4121_),
    .ZN(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4805_ (.A1(_4030_),
    .A2(_4038_),
    .ZN(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4806_ (.A1(_3869_),
    .A2(_4037_),
    .B(_4123_),
    .ZN(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4807_ (.A1(_4054_),
    .A2(_4048_),
    .A3(_4064_),
    .ZN(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4808_ (.A1(_4054_),
    .A2(_4048_),
    .B(_4064_),
    .ZN(_4126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4809_ (.A1(_4053_),
    .A2(_4125_),
    .B(_4126_),
    .ZN(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4810_ (.A1(_3841_),
    .A2(_3844_),
    .ZN(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4811_ (.A1(_4112_),
    .A2(_3604_),
    .ZN(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4812_ (.I(_3293_),
    .Z(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4813_ (.A1(_3849_),
    .A2(_4130_),
    .ZN(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4814_ (.A1(_4128_),
    .A2(_4129_),
    .A3(_4131_),
    .ZN(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4815_ (.I(_3867_),
    .Z(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4816_ (.A1(_3859_),
    .A2(_4133_),
    .ZN(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4817_ (.I(_4034_),
    .ZN(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4818_ (.A1(_3111_),
    .A2(_4135_),
    .ZN(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4819_ (.I(_4135_),
    .Z(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4820_ (.A1(_3872_),
    .A2(_3122_),
    .B1(_4137_),
    .B2(_3859_),
    .ZN(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4821_ (.A1(_4134_),
    .A2(_4136_),
    .B1(_4138_),
    .B2(_4032_),
    .ZN(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4822_ (.A1(_2685_),
    .A2(_3862_),
    .ZN(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4823_ (.A1(_4031_),
    .A2(_3872_),
    .ZN(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4824_ (.A1(_4136_),
    .A2(_4140_),
    .A3(_4141_),
    .ZN(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4825_ (.A1(_4139_),
    .A2(_4142_),
    .Z(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4826_ (.A1(_4132_),
    .A2(_4143_),
    .ZN(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4827_ (.A1(_4127_),
    .A2(_4144_),
    .ZN(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4828_ (.A1(_4124_),
    .A2(_4145_),
    .Z(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4829_ (.A1(_4050_),
    .A2(_4099_),
    .ZN(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4830_ (.A1(_4050_),
    .A2(_4099_),
    .ZN(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4831_ (.A1(_4065_),
    .A2(_4147_),
    .B(_4148_),
    .ZN(_4149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4832_ (.I(_3807_),
    .Z(_4150_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4833_ (.A1(_4057_),
    .A2(_4058_),
    .ZN(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4834_ (.A1(\A[2][7] ),
    .A2(_4078_),
    .B1(_3894_),
    .B2(_4077_),
    .ZN(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4835_ (.A1(_4150_),
    .A2(_4151_),
    .A3(_4152_),
    .B1(_4057_),
    .B2(_4058_),
    .ZN(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4836_ (.A1(_4044_),
    .A2(_4074_),
    .Z(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4837_ (.A1(_4046_),
    .A2(_4068_),
    .ZN(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4838_ (.A1(_4154_),
    .A2(_4082_),
    .B(_4155_),
    .ZN(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4839_ (.I(_4009_),
    .Z(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4840_ (.I(_4066_),
    .Z(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4841_ (.A1(_4158_),
    .A2(_4152_),
    .ZN(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4842_ (.A1(_4157_),
    .A2(_4159_),
    .ZN(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4843_ (.I(_4056_),
    .Z(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4844_ (.A1(_0042_),
    .A2(_4161_),
    .ZN(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4845_ (.A1(_4160_),
    .A2(_4162_),
    .Z(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4846_ (.A1(_4156_),
    .A2(_4163_),
    .Z(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4847_ (.A1(_4153_),
    .A2(_4164_),
    .Z(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4848_ (.A1(_4095_),
    .A2(_4097_),
    .ZN(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4849_ (.A1(_3970_),
    .A2(_3984_),
    .A3(_4166_),
    .B1(_4098_),
    .B2(_4083_),
    .ZN(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4850_ (.I(_3804_),
    .Z(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4851_ (.I(_4168_),
    .Z(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4852_ (.A1(_3917_),
    .A2(_3762_),
    .A3(_4169_),
    .ZN(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4853_ (.A1(_4068_),
    .A2(_4170_),
    .Z(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4854_ (.A1(_3948_),
    .A2(_3936_),
    .ZN(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4855_ (.I(_4172_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4856_ (.I(_4010_),
    .Z(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4857_ (.A1(_0043_),
    .A2(_4173_),
    .ZN(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4858_ (.A1(_4171_),
    .A2(_4174_),
    .Z(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4859_ (.I(_4092_),
    .Z(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4860_ (.A1(_3978_),
    .A2(_4091_),
    .A3(_4176_),
    .ZN(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4861_ (.A1(_4094_),
    .A2(_4097_),
    .B(_4177_),
    .ZN(_4178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4862_ (.I(_4092_),
    .Z(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4863_ (.A1(_3971_),
    .A2(\C[3][8] ),
    .ZN(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _4864_ (.A1(_3948_),
    .A2(_3824_),
    .A3(_4179_),
    .A4(_4180_),
    .Z(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4865_ (.I(_4092_),
    .Z(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4866_ (.A1(_3777_),
    .A2(_3823_),
    .A3(_4182_),
    .B1(_4180_),
    .B2(_4087_),
    .ZN(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4867_ (.A1(_4181_),
    .A2(_4183_),
    .ZN(_4184_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4868_ (.A1(_3793_),
    .A2(_3937_),
    .A3(_3980_),
    .ZN(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4869_ (.A1(_4178_),
    .A2(_4184_),
    .A3(_4185_),
    .Z(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4870_ (.A1(_4175_),
    .A2(_4186_),
    .Z(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4871_ (.A1(_4167_),
    .A2(_4187_),
    .Z(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4872_ (.A1(_4165_),
    .A2(_4188_),
    .Z(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4873_ (.A1(_4146_),
    .A2(_4149_),
    .A3(_4189_),
    .Z(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4874_ (.A1(_4122_),
    .A2(_4190_),
    .Z(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4875_ (.A1(_4120_),
    .A2(_4191_),
    .ZN(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4876_ (.A1(_4105_),
    .A2(_4192_),
    .Z(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4877_ (.A1(_3911_),
    .A2(_4193_),
    .ZN(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4878_ (.I(_2963_),
    .Z(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4879_ (.I(_4195_),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4880_ (.A1(_0059_),
    .A2(_3870_),
    .ZN(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4881_ (.A1(_3144_),
    .A2(_4196_),
    .ZN(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4882_ (.I(_3848_),
    .Z(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4883_ (.A1(_2460_),
    .A2(_4198_),
    .ZN(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4884_ (.I(_2941_),
    .Z(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4885_ (.A1(_3056_),
    .A2(_3089_),
    .B(_3794_),
    .C(_4200_),
    .ZN(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4886_ (.I(_3844_),
    .Z(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4887_ (.A1(_4070_),
    .A2(_4202_),
    .A3(_3856_),
    .A4(_3857_),
    .ZN(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4888_ (.A1(_4201_),
    .A2(_4203_),
    .Z(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4889_ (.A1(_4199_),
    .A2(_4204_),
    .ZN(_4205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4890_ (.A1(_4197_),
    .A2(_4205_),
    .ZN(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4891_ (.I(_3840_),
    .Z(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4892_ (.I(_4207_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4893_ (.A1(_0028_),
    .A2(_3240_),
    .ZN(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4894_ (.A1(_4206_),
    .A2(_4208_),
    .Z(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4895_ (.A1(_4206_),
    .A2(_4208_),
    .Z(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4896_ (.A1(_3510_),
    .A2(_0029_),
    .A3(_4210_),
    .ZN(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4897_ (.A1(_4209_),
    .A2(_4211_),
    .Z(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4898_ (.I(_3956_),
    .Z(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4899_ (.I(_3757_),
    .Z(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4900_ (.I(_4214_),
    .Z(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4901_ (.A1(_4070_),
    .A2(_4213_),
    .A3(_4215_),
    .ZN(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4902_ (.A1(_3774_),
    .A2(_4216_),
    .Z(_4217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4903_ (.I(_4071_),
    .Z(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4904_ (.A1(_4218_),
    .A2(_3809_),
    .ZN(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4905_ (.A1(_3794_),
    .A2(_4002_),
    .A3(_3799_),
    .ZN(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4906_ (.A1(_3791_),
    .A2(_4220_),
    .ZN(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4907_ (.A1(_4217_),
    .A2(_4219_),
    .B(_4221_),
    .ZN(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4908_ (.A1(_3801_),
    .A2(_3810_),
    .Z(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4909_ (.A1(_4222_),
    .A2(_4223_),
    .ZN(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4910_ (.A1(_3865_),
    .A2(_3884_),
    .Z(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4911_ (.A1(_4224_),
    .A2(_4225_),
    .ZN(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4912_ (.I(_3888_),
    .Z(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4913_ (.A1(_4227_),
    .A2(_3905_),
    .ZN(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4914_ (.A1(_4228_),
    .A2(_3662_),
    .ZN(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4915_ (.A1(_4226_),
    .A2(_4229_),
    .ZN(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4916_ (.A1(_4226_),
    .A2(_4229_),
    .ZN(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4917_ (.A1(_4212_),
    .A2(_4230_),
    .B(_4231_),
    .ZN(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4918_ (.A1(_4212_),
    .A2(_4230_),
    .Z(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4919_ (.I(_4233_),
    .ZN(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4920_ (.A1(_4224_),
    .A2(_4225_),
    .Z(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4921_ (.I(_4235_),
    .ZN(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4922_ (.A1(_4222_),
    .A2(_4223_),
    .ZN(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4923_ (.A1(_3997_),
    .A2(_3818_),
    .ZN(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4924_ (.I(_3928_),
    .Z(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4925_ (.A1(\C[3][3] ),
    .A2(_4239_),
    .ZN(_4240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4926_ (.A1(_4238_),
    .A2(_4240_),
    .ZN(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4927_ (.I(_3927_),
    .Z(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4928_ (.A1(\C[3][4] ),
    .A2(_4242_),
    .ZN(_4243_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4929_ (.A1(_3918_),
    .A2(_3923_),
    .A3(_4243_),
    .ZN(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4930_ (.A1(_4241_),
    .A2(_4244_),
    .Z(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4931_ (.I(_4245_),
    .ZN(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4932_ (.A1(_4241_),
    .A2(_4244_),
    .ZN(_4247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4933_ (.A1(_4237_),
    .A2(_4246_),
    .B(_4247_),
    .ZN(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4934_ (.A1(_3930_),
    .A2(_3941_),
    .A3(_3914_),
    .ZN(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4935_ (.A1(_4248_),
    .A2(_4249_),
    .ZN(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4936_ (.A1(_4248_),
    .A2(_4249_),
    .ZN(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4937_ (.A1(_4236_),
    .A2(_4250_),
    .B(_4251_),
    .ZN(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4938_ (.A1(_3944_),
    .A2(_4019_),
    .A3(_3913_),
    .ZN(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4939_ (.A1(_4252_),
    .A2(_4253_),
    .ZN(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4940_ (.A1(_4252_),
    .A2(_4253_),
    .ZN(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4941_ (.A1(_4234_),
    .A2(_4254_),
    .B(_4255_),
    .ZN(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4942_ (.A1(_3912_),
    .A2(_4103_),
    .Z(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4943_ (.A1(_4256_),
    .A2(_4257_),
    .Z(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4944_ (.A1(_4256_),
    .A2(_4257_),
    .Z(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4945_ (.A1(_4232_),
    .A2(_4258_),
    .B(_4259_),
    .ZN(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4946_ (.A1(_4194_),
    .A2(_4260_),
    .Z(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4947_ (.I(_3845_),
    .Z(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4948_ (.I(_4262_),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4949_ (.A1(_0027_),
    .A2(_3240_),
    .ZN(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4950_ (.A1(_0058_),
    .A2(_3871_),
    .A3(_4201_),
    .ZN(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4951_ (.A1(_4263_),
    .A2(_4264_),
    .ZN(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4952_ (.A1(_4263_),
    .A2(_4264_),
    .ZN(_4266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4953_ (.A1(_0028_),
    .A2(_3889_),
    .ZN(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4954_ (.A1(_4266_),
    .A2(_4267_),
    .ZN(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4955_ (.A1(_4265_),
    .A2(_4268_),
    .ZN(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4956_ (.A1(_3762_),
    .A2(_3922_),
    .A3(_3767_),
    .ZN(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4957_ (.A1(_3814_),
    .A2(_4007_),
    .ZN(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4958_ (.A1(_4270_),
    .A2(_4271_),
    .Z(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4959_ (.I(_3953_),
    .Z(_4273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4960_ (.A1(_3809_),
    .A2(_4273_),
    .ZN(_4274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4961_ (.I(_3965_),
    .Z(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4962_ (.A1(_4275_),
    .A2(_4215_),
    .A3(_4220_),
    .ZN(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4963_ (.A1(_4272_),
    .A2(_4274_),
    .B(_4276_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4964_ (.A1(_3791_),
    .A2(_4220_),
    .B1(_4216_),
    .B2(_3774_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4965_ (.A1(_0150_),
    .A2(_4219_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4966_ (.A1(_0149_),
    .A2(_0151_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4967_ (.A1(_4199_),
    .A2(_4204_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4968_ (.A1(_0152_),
    .A2(_0153_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4969_ (.A1(_4227_),
    .A2(_3326_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4970_ (.A1(_0155_),
    .A2(_4210_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4971_ (.A1(_0154_),
    .A2(_0156_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4972_ (.A1(_0154_),
    .A2(_0156_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4973_ (.A1(_4269_),
    .A2(_0157_),
    .B(_0158_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4974_ (.A1(_0154_),
    .A2(_0156_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4975_ (.A1(_4269_),
    .A2(_0160_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4976_ (.A1(_0152_),
    .A2(_0153_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4977_ (.A1(_0149_),
    .A2(_0151_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4978_ (.A1(_4238_),
    .A2(_4240_),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4979_ (.A1(_4222_),
    .A2(_4223_),
    .A3(_4245_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4980_ (.A1(_0163_),
    .A2(_0164_),
    .B(_0165_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4981_ (.A1(_0163_),
    .A2(_0164_),
    .A3(_0165_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4982_ (.A1(_0162_),
    .A2(_0166_),
    .B(_0167_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4983_ (.A1(_4248_),
    .A2(_4249_),
    .A3(_4235_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4984_ (.A1(_0168_),
    .A2(_0169_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4985_ (.A1(_0168_),
    .A2(_0169_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4986_ (.A1(_0161_),
    .A2(_0170_),
    .B(_0171_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4987_ (.A1(_4252_),
    .A2(_4253_),
    .A3(_4233_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4988_ (.A1(_0172_),
    .A2(_0173_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4989_ (.A1(_0172_),
    .A2(_0173_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4990_ (.A1(_0159_),
    .A2(_0174_),
    .B(_0175_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4991_ (.A1(_4232_),
    .A2(_4258_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4992_ (.A1(_0176_),
    .A2(_0177_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4993_ (.A1(\B[1][0] ),
    .A2(_3764_),
    .B1(_3391_),
    .B2(_3765_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4994_ (.A1(_3979_),
    .A2(_0179_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4995_ (.I(_4002_),
    .Z(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4996_ (.A1(_3979_),
    .A2(_3799_),
    .B1(_4150_),
    .B2(_0181_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4997_ (.A1(_4270_),
    .A2(_0180_),
    .B(_0182_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4998_ (.I(_4242_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4999_ (.I(_0184_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5000_ (.I(_0185_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5001_ (.A1(\C[3][1] ),
    .A2(_0186_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5002_ (.A1(_0183_),
    .A2(_0187_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5003_ (.A1(\C[3][0] ),
    .A2(_0186_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5004_ (.A1(_0180_),
    .A2(_0189_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5005_ (.A1(_0188_),
    .A2(_0190_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5006_ (.A1(_0058_),
    .A2(_3882_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5007_ (.A1(_4270_),
    .A2(_4271_),
    .A3(_4274_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5008_ (.A1(_4270_),
    .A2(_0180_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5009_ (.A1(\C[3][2] ),
    .A2(_0184_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5010_ (.A1(_0193_),
    .A2(_0194_),
    .A3(_0195_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5011_ (.A1(_0183_),
    .A2(_0187_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5012_ (.A1(_0192_),
    .A2(_0196_),
    .A3(_0197_),
    .Z(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5013_ (.I(_3133_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5014_ (.I(_0199_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5015_ (.I(_0200_),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5016_ (.I(_0201_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5017_ (.I(_3904_),
    .Z(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5018_ (.I(_2889_),
    .Z(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5019_ (.A1(_0203_),
    .A2(_4227_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5020_ (.I(_0204_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5021_ (.I(_4033_),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5022_ (.I(_0206_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5023_ (.I(_3488_),
    .Z(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5024_ (.A1(_0207_),
    .A2(_0208_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5025_ (.A1(_0025_),
    .A2(_0202_),
    .A3(_0205_),
    .A4(_0209_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5026_ (.I(_3904_),
    .Z(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5027_ (.A1(_0201_),
    .A2(_0211_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5028_ (.A1(_0205_),
    .A2(_0212_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5029_ (.I(_0203_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5030_ (.I(_0025_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5031_ (.A1(_0214_),
    .A2(_0208_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5032_ (.A1(_0026_),
    .A2(_0207_),
    .A3(_4117_),
    .A4(_0215_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5033_ (.A1(_0210_),
    .A2(_0213_),
    .A3(_0216_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5034_ (.A1(_0191_),
    .A2(_0198_),
    .A3(_0217_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5035_ (.A1(_0188_),
    .A2(_0190_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5036_ (.I(_3882_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5037_ (.I(_3903_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5038_ (.A1(_0024_),
    .A2(_0220_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5039_ (.A1(_0215_),
    .A2(_0221_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5040_ (.A1(_0219_),
    .A2(_0222_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5041_ (.A1(_0180_),
    .A2(_0189_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5042_ (.A1(_0209_),
    .A2(_0224_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5043_ (.A1(_0223_),
    .A2(_0225_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5044_ (.A1(_0218_),
    .A2(_0226_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5045_ (.I(_0227_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5046_ (.I(_0222_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5047_ (.A1(_0219_),
    .A2(_0229_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5048_ (.A1(_0218_),
    .A2(_0230_),
    .Z(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5049_ (.A1(_0191_),
    .A2(_0198_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5050_ (.A1(_0191_),
    .A2(_0198_),
    .Z(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5051_ (.A1(_0217_),
    .A2(_0232_),
    .B(_0233_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5052_ (.A1(_0196_),
    .A2(_0197_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5053_ (.A1(_0196_),
    .A2(_0197_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5054_ (.A1(_0192_),
    .A2(_0235_),
    .B(_0236_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5055_ (.A1(_0149_),
    .A2(_0151_),
    .A3(_0164_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5056_ (.A1(_0193_),
    .A2(_0194_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5057_ (.A1(_0193_),
    .A2(_0194_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5058_ (.A1(_0239_),
    .A2(_0240_),
    .A3(_0195_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5059_ (.A1(_4113_),
    .A2(_0200_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5060_ (.A1(_4196_),
    .A2(_0242_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5061_ (.A1(_0239_),
    .A2(_0243_),
    .Z(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5062_ (.A1(_0238_),
    .A2(_0241_),
    .A3(_0244_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5063_ (.A1(_4263_),
    .A2(_0204_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5064_ (.A1(_0205_),
    .A2(_0246_),
    .A3(_0212_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5065_ (.I(_0247_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5066_ (.A1(_0027_),
    .A2(_0056_),
    .B1(_0220_),
    .B2(_0026_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5067_ (.A1(_0025_),
    .A2(_4117_),
    .B(_4263_),
    .C(_0205_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5068_ (.A1(_0248_),
    .A2(_0249_),
    .A3(_0250_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5069_ (.A1(_0237_),
    .A2(_0245_),
    .A3(_0251_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5070_ (.A1(_0210_),
    .A2(_0234_),
    .A3(_0252_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5071_ (.A1(_0231_),
    .A2(_0253_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5072_ (.A1(_0231_),
    .A2(_0253_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5073_ (.A1(_0228_),
    .A2(_0254_),
    .B(_0255_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5074_ (.A1(_0234_),
    .A2(_0252_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5075_ (.A1(_0234_),
    .A2(_0252_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5076_ (.A1(_0210_),
    .A2(_0257_),
    .B(_0258_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5077_ (.I(_0251_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5078_ (.A1(_0237_),
    .A2(_0245_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5079_ (.A1(_0237_),
    .A2(_0245_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5080_ (.A1(_0260_),
    .A2(_0261_),
    .B(_0262_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5081_ (.I(_0244_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5082_ (.A1(_0238_),
    .A2(_0241_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5083_ (.A1(_0238_),
    .A2(_0241_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5084_ (.A1(_0264_),
    .A2(_0265_),
    .B(_0266_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5085_ (.A1(_0163_),
    .A2(_0164_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5086_ (.A1(_0268_),
    .A2(_0165_),
    .A3(_0162_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5087_ (.A1(_0239_),
    .A2(_0243_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5088_ (.A1(_4266_),
    .A2(_4267_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5089_ (.A1(_0270_),
    .A2(_0271_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5090_ (.A1(_0246_),
    .A2(_0272_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5091_ (.A1(_0267_),
    .A2(_0269_),
    .A3(_0273_),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5092_ (.A1(_0248_),
    .A2(_0263_),
    .A3(_0274_),
    .Z(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5093_ (.A1(_0259_),
    .A2(_0275_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5094_ (.A1(_0259_),
    .A2(_0275_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5095_ (.A1(_0256_),
    .A2(_0276_),
    .B(_0277_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5096_ (.A1(_0263_),
    .A2(_0274_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5097_ (.A1(_0263_),
    .A2(_0274_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5098_ (.A1(_0247_),
    .A2(_0279_),
    .B(_0280_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5099_ (.I(_0273_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5100_ (.A1(_0267_),
    .A2(_0269_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5101_ (.A1(_0267_),
    .A2(_0269_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5102_ (.A1(_0282_),
    .A2(_0283_),
    .B(_0284_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5103_ (.A1(_0161_),
    .A2(_0170_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5104_ (.A1(_0270_),
    .A2(_0271_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5105_ (.A1(_0246_),
    .A2(_0272_),
    .B(_0287_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5106_ (.I(_0288_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5107_ (.A1(_0285_),
    .A2(_0286_),
    .A3(_0289_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5108_ (.A1(_0281_),
    .A2(_0290_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5109_ (.A1(_0281_),
    .A2(_0290_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5110_ (.A1(_0278_),
    .A2(_0291_),
    .B(_0292_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5111_ (.A1(_0285_),
    .A2(_0286_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5112_ (.A1(_0285_),
    .A2(_0286_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5113_ (.A1(_0289_),
    .A2(_0294_),
    .B(_0295_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5114_ (.A1(_0159_),
    .A2(_0174_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5115_ (.A1(_0296_),
    .A2(_0297_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5116_ (.A1(_0296_),
    .A2(_0297_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5117_ (.A1(_0176_),
    .A2(_0177_),
    .B1(_0293_),
    .B2(_0298_),
    .C(_0299_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5118_ (.A1(_0178_),
    .A2(_0300_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5119_ (.A1(_4261_),
    .A2(_0301_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5120_ (.I(_0302_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5121_ (.A1(_3727_),
    .A2(_2276_),
    .A3(_2556_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5122_ (.I(_0303_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5123_ (.A1(_2233_),
    .A2(_2254_),
    .A3(_3747_),
    .A4(_2287_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5124_ (.I(_0305_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5125_ (.A1(_3271_),
    .A2(_0304_),
    .B1(_0306_),
    .B2(\B[2][5] ),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5126_ (.I(_0307_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5127_ (.A1(_4033_),
    .A2(_0308_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5128_ (.I(_4031_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5129_ (.I(_0303_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5130_ (.I(_0305_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5131_ (.A1(_2599_),
    .A2(net45),
    .B1(_0312_),
    .B2(\B[2][3] ),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5132_ (.I(_0313_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5133_ (.I(_0314_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5134_ (.A1(_0310_),
    .A2(_0315_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5135_ (.A1(_3819_),
    .A2(net45),
    .B1(_0312_),
    .B2(\B[2][4] ),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5136_ (.I(_0317_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5137_ (.I(_0318_),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5138_ (.I(_0319_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5139_ (.A1(_3875_),
    .A2(_0320_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5140_ (.A1(_0316_),
    .A2(_0321_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5141_ (.A1(_0316_),
    .A2(_0321_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5142_ (.A1(_0309_),
    .A2(_0322_),
    .B(_0323_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5143_ (.A1(net44),
    .A2(_0304_),
    .B1(_0306_),
    .B2(\B[2][6] ),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5144_ (.I(_0325_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5145_ (.I(_0326_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5146_ (.A1(_0206_),
    .A2(_0326_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5147_ (.A1(_0324_),
    .A2(_0328_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _5148_ (.A1(_2610_),
    .A2(_2265_),
    .Z(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5149_ (.I(_0330_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5150_ (.A1(_3982_),
    .A2(_3892_),
    .A3(_0331_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5151_ (.A1(_3892_),
    .A2(_3391_),
    .A3(_0331_),
    .B1(_0332_),
    .B2(\B[0][0] ),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5152_ (.I(_0333_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5153_ (.I(_3778_),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5154_ (.I(_0335_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5155_ (.A1(\A[2][6] ),
    .A2(_4078_),
    .B1(net44),
    .B2(_4077_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5156_ (.A1(_0336_),
    .A2(_0337_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5157_ (.I(_0338_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5158_ (.I(_0022_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _5159_ (.A1(_0207_),
    .A2(_0324_),
    .A3(_0327_),
    .B1(_0329_),
    .B2(_0334_),
    .B3(_0339_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5160_ (.A1(_0309_),
    .A2(_0322_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5161_ (.I(_0310_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5162_ (.A1(_2816_),
    .A2(_0311_),
    .B1(_0312_),
    .B2(\B[2][2] ),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5163_ (.I(_0343_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5164_ (.I(_0344_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5165_ (.I(_0330_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _5166_ (.A1(_2492_),
    .A2(_3782_),
    .A3(_0346_),
    .B(\B[0][2] ),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5167_ (.I(_0347_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5168_ (.A1(_2610_),
    .A2(_2362_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5169_ (.I(_0349_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5170_ (.A1(_3456_),
    .A2(_2816_),
    .A3(_0350_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5171_ (.I(_0351_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5172_ (.A1(_0348_),
    .A2(_0352_),
    .B(_3593_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5173_ (.I(_0353_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5174_ (.I(_0354_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5175_ (.I(_3773_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5176_ (.A1(_0342_),
    .A2(_0345_),
    .B1(_0355_),
    .B2(_0356_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _5177_ (.A1(_3853_),
    .A2(_2578_),
    .A3(_0346_),
    .B(\B[0][1] ),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5178_ (.A1(_3456_),
    .A2(_3078_),
    .A3(_0350_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5179_ (.A1(_0358_),
    .A2(_0359_),
    .B(_3990_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5180_ (.A1(_4072_),
    .A2(_0360_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5181_ (.I(_0344_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5182_ (.I(_0362_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5183_ (.I(_0363_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5184_ (.A1(_0356_),
    .A2(_3848_),
    .A3(_0364_),
    .A4(_0355_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5185_ (.A1(_0357_),
    .A2(_0361_),
    .B(_0365_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5186_ (.A1(_3845_),
    .A2(_0362_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5187_ (.A1(_4071_),
    .A2(_0354_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5188_ (.A1(_4169_),
    .A2(_0360_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5189_ (.A1(_0367_),
    .A2(_0368_),
    .A3(_0369_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5190_ (.A1(_0366_),
    .A2(_0370_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5191_ (.A1(_0366_),
    .A2(_0370_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5192_ (.A1(_0341_),
    .A2(_0371_),
    .B(_0372_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5193_ (.I(_2706_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5194_ (.A1(_3797_),
    .A2(_0311_),
    .B1(_0312_),
    .B2(\B[2][1] ),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _5195_ (.I(_0375_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5196_ (.I(_0376_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5197_ (.I(_0377_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _5198_ (.A1(_3853_),
    .A2(_2578_),
    .A3(_0346_),
    .B(\B[0][4] ),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5199_ (.I(_0349_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _5200_ (.A1(_3048_),
    .A2(_2982_),
    .A3(_0380_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5201_ (.A1(_0379_),
    .A2(_0381_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5202_ (.I(_0382_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5203_ (.I(_0383_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5204_ (.A1(_0374_),
    .A2(_0378_),
    .B1(_0384_),
    .B2(_3997_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5205_ (.I(_3956_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _5206_ (.A1(_3531_),
    .A2(_2786_),
    .A3(_0330_),
    .B(\B[0][3] ),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5207_ (.A1(_2513_),
    .A2(_2599_),
    .A3(_0350_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5208_ (.A1(_0387_),
    .A2(_0388_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5209_ (.A1(_3701_),
    .A2(_0389_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _5210_ (.I(_0390_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5211_ (.I(_0391_),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5212_ (.I(_0392_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5213_ (.A1(_0386_),
    .A2(_0393_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5214_ (.A1(_4275_),
    .A2(_0374_),
    .A3(_0377_),
    .A4(_0384_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5215_ (.A1(_0385_),
    .A2(_0394_),
    .B(_0395_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5216_ (.I(_3840_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5217_ (.I(_0397_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5218_ (.A1(_0398_),
    .A2(_0377_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _5219_ (.A1(_0379_),
    .A2(_0381_),
    .B(_3946_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5220_ (.I(_0400_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5221_ (.A1(_4213_),
    .A2(_0401_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5222_ (.I(_0391_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5223_ (.A1(_0356_),
    .A2(_0403_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5224_ (.A1(_0399_),
    .A2(_0402_),
    .A3(_0404_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5225_ (.A1(_0396_),
    .A2(_0405_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5226_ (.A1(_3848_),
    .A2(_0320_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5227_ (.I(_0307_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5228_ (.I(_0408_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5229_ (.A1(_3133_),
    .A2(_0409_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5230_ (.A1(_2717_),
    .A2(_0315_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5231_ (.A1(_0407_),
    .A2(_0410_),
    .A3(_0411_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5232_ (.I(_0362_),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5233_ (.I(_0413_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5234_ (.I(_0353_),
    .Z(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5235_ (.I(_0415_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5236_ (.A1(_4262_),
    .A2(_0414_),
    .B1(_0034_),
    .B2(_4073_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5237_ (.A1(_4073_),
    .A2(_4262_),
    .A3(_0414_),
    .A4(_0034_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5238_ (.A1(_0416_),
    .A2(_0369_),
    .B(_0417_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5239_ (.I(_3841_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5240_ (.A1(_0419_),
    .A2(_0414_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5241_ (.A1(_3806_),
    .A2(_0415_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5242_ (.I(_3831_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5243_ (.I(_0360_),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5244_ (.A1(_0422_),
    .A2(_0423_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5245_ (.A1(_0420_),
    .A2(_0421_),
    .A3(_0424_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5246_ (.A1(_0412_),
    .A2(_0418_),
    .A3(_0425_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5247_ (.A1(_0406_),
    .A2(_0426_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5248_ (.A1(_0406_),
    .A2(_0426_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5249_ (.A1(_0373_),
    .A2(_0427_),
    .B(_0428_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5250_ (.I(_4159_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5251_ (.A1(_3890_),
    .A2(net5),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5252_ (.A1(_3892_),
    .A2(_0331_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5253_ (.A1(_3413_),
    .A2(_3467_),
    .A3(_0380_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5254_ (.I(\B[0][0] ),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5255_ (.A1(_0430_),
    .A2(_0431_),
    .B1(_0432_),
    .B2(_0433_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5256_ (.I(_0434_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5257_ (.I(_0435_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5258_ (.A1(_0023_),
    .A2(_0436_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5259_ (.I(_0315_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5260_ (.A1(_4262_),
    .A2(_0051_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5261_ (.A1(_0407_),
    .A2(_0438_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5262_ (.A1(_2695_),
    .A2(_0319_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5263_ (.A1(_0316_),
    .A2(_0440_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5264_ (.A1(_0410_),
    .A2(_0439_),
    .B(_0441_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5265_ (.I(_0325_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5266_ (.I(_0443_),
    .Z(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5267_ (.I(_0444_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5268_ (.A1(_0201_),
    .A2(_0445_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5269_ (.A1(_0442_),
    .A2(_0446_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5270_ (.A1(_0437_),
    .A2(_0447_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5271_ (.A1(_0429_),
    .A2(_0448_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5272_ (.A1(_0429_),
    .A2(_0448_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5273_ (.A1(_0340_),
    .A2(_0449_),
    .B(_0450_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5274_ (.A1(_0340_),
    .A2(_0449_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5275_ (.I(_0452_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5276_ (.A1(_0406_),
    .A2(_0373_),
    .A3(_0426_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5277_ (.A1(_0396_),
    .A2(_0405_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5278_ (.I(_4089_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5279_ (.I(_0456_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5280_ (.A1(_0457_),
    .A2(\C[2][3] ),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5281_ (.I(\B[2][0] ),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5282_ (.A1(_0430_),
    .A2(_0304_),
    .B1(_0306_),
    .B2(_0459_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5283_ (.I(_0460_),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5284_ (.I(_0461_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5285_ (.A1(_0374_),
    .A2(_0458_),
    .A3(_0462_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5286_ (.A1(_3983_),
    .A2(\C[2][4] ),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5287_ (.A1(_0398_),
    .A2(_0461_),
    .A3(_0464_),
    .Z(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5288_ (.I(_0460_),
    .Z(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5289_ (.I(_0466_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5290_ (.I(_3975_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5291_ (.I(_0468_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5292_ (.A1(_4207_),
    .A2(_0467_),
    .B1(_0464_),
    .B2(_0469_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5293_ (.A1(_0463_),
    .A2(_0465_),
    .A3(_0470_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5294_ (.I(_0460_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5295_ (.I(_4089_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5296_ (.A1(_0473_),
    .A2(\C[2][5] ),
    .Z(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5297_ (.A1(_3304_),
    .A2(_0472_),
    .A3(_0474_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5298_ (.I(_3974_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5299_ (.A1(_4130_),
    .A2(_0472_),
    .B1(_0474_),
    .B2(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5300_ (.A1(_0475_),
    .A2(_0477_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _5301_ (.A1(_3531_),
    .A2(_2786_),
    .A3(_0330_),
    .B(\B[0][5] ),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5302_ (.A1(_3456_),
    .A2(_3260_),
    .A3(_0350_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5303_ (.A1(_0479_),
    .A2(_0480_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5304_ (.A1(_3997_),
    .A2(_0481_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5305_ (.A1(_0465_),
    .A2(_0478_),
    .A3(_0482_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5306_ (.A1(_0471_),
    .A2(_0483_),
    .Z(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5307_ (.A1(_0471_),
    .A2(_0483_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5308_ (.A1(_0455_),
    .A2(_0484_),
    .B(_0485_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5309_ (.I(_0400_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5310_ (.I(_0487_),
    .Z(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5311_ (.I(_0488_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5312_ (.I(_3922_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5313_ (.A1(_4207_),
    .A2(_0378_),
    .B1(_0036_),
    .B2(_0489_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5314_ (.A1(_0489_),
    .A2(_4207_),
    .A3(_0378_),
    .A4(_0036_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5315_ (.A1(_0490_),
    .A2(_0404_),
    .B(_0491_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5316_ (.I(_0376_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5317_ (.A1(_3315_),
    .A2(_0493_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5318_ (.A1(_3773_),
    .A2(_0401_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5319_ (.A1(_4072_),
    .A2(_0393_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5320_ (.A1(_0494_),
    .A2(_0495_),
    .A3(_0496_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5321_ (.I(_0461_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5322_ (.A1(_0419_),
    .A2(_0498_),
    .A3(_0464_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5323_ (.A1(_0475_),
    .A2(_0477_),
    .B(_0499_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5324_ (.A1(_0499_),
    .A2(_0475_),
    .A3(_0477_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5325_ (.A1(_0500_),
    .A2(_0482_),
    .B(_0501_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5326_ (.A1(_3315_),
    .A2(_0461_),
    .A3(_0474_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5327_ (.A1(_3542_),
    .A2(_2794_),
    .A3(_0331_),
    .B(\B[0][6] ),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5328_ (.A1(_2755_),
    .A2(_3562_),
    .A3(_0380_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5329_ (.A1(_0504_),
    .A2(_0505_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5330_ (.A1(_3813_),
    .A2(_0506_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5331_ (.A1(_0479_),
    .A2(_0480_),
    .B(_3990_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5332_ (.I(_0508_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5333_ (.A1(_3921_),
    .A2(_0509_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5334_ (.A1(_0507_),
    .A2(_0510_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5335_ (.I(net37),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5336_ (.I(_3854_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5337_ (.I(_0513_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5338_ (.A1(_0514_),
    .A2(\C[2][6] ),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _5339_ (.A1(_0512_),
    .A2(_0472_),
    .A3(_0515_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5340_ (.A1(_0512_),
    .A2(_0466_),
    .B1(_0515_),
    .B2(_3976_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5341_ (.A1(_0516_),
    .A2(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5342_ (.A1(_0503_),
    .A2(_0511_),
    .A3(_0518_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5343_ (.A1(_0502_),
    .A2(_0519_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5344_ (.A1(_0492_),
    .A2(_0497_),
    .A3(_0520_),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5345_ (.A1(_0486_),
    .A2(_0521_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5346_ (.A1(_0486_),
    .A2(_0521_),
    .Z(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5347_ (.A1(_0454_),
    .A2(_0522_),
    .B(_0523_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5348_ (.A1(_0418_),
    .A2(_0425_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5349_ (.A1(_0418_),
    .A2(_0425_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5350_ (.A1(_0412_),
    .A2(_0525_),
    .B(_0526_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5351_ (.A1(_0492_),
    .A2(_0497_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5352_ (.I(_0314_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5353_ (.A1(_0397_),
    .A2(_0529_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5354_ (.A1(_0310_),
    .A2(_0408_),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5355_ (.A1(_0440_),
    .A2(_0530_),
    .A3(_0531_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5356_ (.I(_0353_),
    .Z(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5357_ (.A1(_3842_),
    .A2(_0413_),
    .B1(_0533_),
    .B2(_4169_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5358_ (.A1(_3806_),
    .A2(_0398_),
    .A3(_0413_),
    .A4(_0533_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5359_ (.A1(_0534_),
    .A2(_0424_),
    .B(_0535_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5360_ (.I(_0362_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5361_ (.A1(_4130_),
    .A2(_0537_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5362_ (.I(_0353_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5363_ (.A1(_4010_),
    .A2(_0539_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5364_ (.I(_4056_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5365_ (.A1(_0541_),
    .A2(_0423_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5366_ (.A1(_0538_),
    .A2(_0540_),
    .A3(_0542_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5367_ (.A1(_0532_),
    .A2(_0536_),
    .A3(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5368_ (.A1(_0528_),
    .A2(_0544_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5369_ (.A1(_0527_),
    .A2(_0545_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5370_ (.A1(_0492_),
    .A2(_0497_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5371_ (.A1(_0528_),
    .A2(_0547_),
    .A3(_0520_),
    .B1(_0519_),
    .B2(_0502_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5372_ (.A1(_0494_),
    .A2(_0495_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5373_ (.I(_0496_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5374_ (.A1(_0494_),
    .A2(_0495_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5375_ (.A1(_0549_),
    .A2(_0550_),
    .B(_0551_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5376_ (.A1(_0507_),
    .A2(_0510_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5377_ (.A1(_3604_),
    .A2(_0376_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5378_ (.A1(_3751_),
    .A2(_0400_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5379_ (.A1(_4168_),
    .A2(_0392_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5380_ (.A1(_0554_),
    .A2(_0555_),
    .A3(_0556_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5381_ (.A1(_0553_),
    .A2(_0557_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5382_ (.A1(_0552_),
    .A2(_0558_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5383_ (.I(_0516_),
    .Z(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5384_ (.A1(_0560_),
    .A2(_0517_),
    .B(_0503_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5385_ (.A1(_0503_),
    .A2(_0560_),
    .A3(_0517_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5386_ (.A1(_0511_),
    .A2(_0561_),
    .B(_0562_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _5387_ (.A1(_3853_),
    .A2(_2578_),
    .A3(_0346_),
    .B(\B[0][7] ),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _5388_ (.A1(_2755_),
    .A2(_3893_),
    .A3(_0380_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5389_ (.A1(_0564_),
    .A2(_0565_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5390_ (.A1(_3978_),
    .A2(_0566_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5391_ (.A1(_0504_),
    .A2(_0505_),
    .B(_3593_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5392_ (.I(_0568_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5393_ (.A1(_3921_),
    .A2(_0569_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5394_ (.I(_0509_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5395_ (.A1(_3953_),
    .A2(_0571_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5396_ (.A1(_0567_),
    .A2(_0570_),
    .A3(_0572_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5397_ (.I(_3896_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5398_ (.A1(_0574_),
    .A2(_0472_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _5399_ (.A1(_3894_),
    .A2(_0304_),
    .B1(_0306_),
    .B2(\B[2][7] ),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5400_ (.I(_0576_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5401_ (.A1(_4033_),
    .A2(_0577_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5402_ (.A1(\C[2][7] ),
    .A2(_4242_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5403_ (.A1(_0575_),
    .A2(_0578_),
    .A3(_0579_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5404_ (.A1(_0516_),
    .A2(_0573_),
    .A3(_0580_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5405_ (.A1(_0559_),
    .A2(_0563_),
    .A3(_0581_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5406_ (.A1(_0548_),
    .A2(_0582_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5407_ (.A1(_0546_),
    .A2(_0583_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5408_ (.A1(_0524_),
    .A2(_0584_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5409_ (.A1(_0524_),
    .A2(_0584_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5410_ (.A1(_0453_),
    .A2(_0585_),
    .B(_0586_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _5411_ (.A1(_0214_),
    .A2(_0327_),
    .A3(_0442_),
    .B1(_0447_),
    .B2(_0437_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5412_ (.A1(_0026_),
    .A2(_0445_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5413_ (.A1(_0398_),
    .A2(_0320_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5414_ (.I(_0590_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5415_ (.A1(_0440_),
    .A2(_0530_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5416_ (.A1(_0411_),
    .A2(_0591_),
    .B1(_0592_),
    .B2(_0531_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5417_ (.A1(_0589_),
    .A2(_0593_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5418_ (.A1(_0528_),
    .A2(_0544_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5419_ (.A1(_0527_),
    .A2(_0545_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5420_ (.A1(_0595_),
    .A2(_0596_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5421_ (.A1(_0594_),
    .A2(_0597_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5422_ (.A1(_0588_),
    .A2(_0598_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5423_ (.A1(_0548_),
    .A2(_0582_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5424_ (.A1(_0546_),
    .A2(_0583_),
    .B(_0600_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5425_ (.A1(_0536_),
    .A2(_0543_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5426_ (.A1(_0536_),
    .A2(_0543_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5427_ (.A1(_0532_),
    .A2(_0602_),
    .B(_0603_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5428_ (.A1(_0507_),
    .A2(_0510_),
    .A3(_0557_),
    .Z(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5429_ (.A1(_0552_),
    .A2(_0558_),
    .B(_0605_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5430_ (.I(_0408_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5431_ (.A1(_2717_),
    .A2(_0607_),
    .Z(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5432_ (.A1(_4130_),
    .A2(_0529_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5433_ (.A1(_0590_),
    .A2(_0609_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5434_ (.A1(_0608_),
    .A2(_0610_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5435_ (.A1(_4026_),
    .A2(_0364_),
    .B1(_0355_),
    .B2(_0422_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5436_ (.A1(_4173_),
    .A2(_4026_),
    .A3(_0364_),
    .A4(_0355_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5437_ (.A1(_0612_),
    .A2(_0542_),
    .B(_0613_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5438_ (.A1(_3615_),
    .A2(_0363_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5439_ (.A1(_4056_),
    .A2(_0354_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5440_ (.A1(_4061_),
    .A2(_0423_),
    .ZN(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5441_ (.A1(_0615_),
    .A2(_0616_),
    .A3(_0617_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5442_ (.A1(_0614_),
    .A2(_0618_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5443_ (.A1(_0611_),
    .A2(_0619_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5444_ (.A1(_0606_),
    .A2(_0620_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5445_ (.A1(_0604_),
    .A2(_0621_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5446_ (.A1(_0563_),
    .A2(_0581_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5447_ (.A1(_0563_),
    .A2(_0581_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5448_ (.A1(_0559_),
    .A2(_0623_),
    .B(_0624_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5449_ (.A1(_0554_),
    .A2(_0555_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5450_ (.A1(_4080_),
    .A2(_0390_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5451_ (.A1(_0554_),
    .A2(_0555_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5452_ (.A1(_0626_),
    .A2(_0627_),
    .B(_0628_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5453_ (.A1(_0564_),
    .A2(_0565_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5454_ (.I(_0630_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5455_ (.I(_0631_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5456_ (.I(_0568_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5457_ (.A1(_3965_),
    .A2(_0632_),
    .B1(_0633_),
    .B2(_4213_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5458_ (.A1(_3965_),
    .A2(_4213_),
    .A3(_0632_),
    .A4(_0633_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5459_ (.A1(_0634_),
    .A2(_0572_),
    .B(_0635_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5460_ (.A1(_0574_),
    .A2(_0493_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5461_ (.A1(_3805_),
    .A2(_0487_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5462_ (.A1(_0422_),
    .A2(_0393_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5463_ (.A1(_0637_),
    .A2(_0638_),
    .A3(_0639_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5464_ (.A1(_0629_),
    .A2(_0636_),
    .A3(_0640_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5465_ (.I(_0573_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5466_ (.A1(_0560_),
    .A2(_0580_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5467_ (.A1(_0560_),
    .A2(_0580_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5468_ (.A1(_0642_),
    .A2(_0643_),
    .B(_0644_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5469_ (.I(_0568_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5470_ (.I(_0646_),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5471_ (.A1(_0564_),
    .A2(_0565_),
    .B(_3946_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5472_ (.I(_0648_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5473_ (.A1(_0386_),
    .A2(_4273_),
    .A3(_0647_),
    .A4(_0649_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5474_ (.I(_0648_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5475_ (.A1(_3772_),
    .A2(_0569_),
    .B1(_0651_),
    .B2(_3956_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5476_ (.A1(_0650_),
    .A2(_0652_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5477_ (.A1(_4071_),
    .A2(_0571_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5478_ (.A1(_0653_),
    .A2(_0654_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5479_ (.I(_0576_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5480_ (.I(_0656_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5481_ (.I(_0657_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5482_ (.A1(\C[2][7] ),
    .A2(_4242_),
    .B1(_0658_),
    .B2(_3860_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5483_ (.A1(\C[2][7] ),
    .A2(_3860_),
    .A3(_3928_),
    .A4(_0658_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5484_ (.A1(_0575_),
    .A2(_0659_),
    .B(_0660_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5485_ (.A1(_3972_),
    .A2(\C[2][8] ),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5486_ (.A1(_3133_),
    .A2(_0657_),
    .A3(_0662_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5487_ (.A1(_3875_),
    .A2(_0658_),
    .B1(_0662_),
    .B2(_0468_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5488_ (.A1(_0663_),
    .A2(_0664_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5489_ (.A1(_0661_),
    .A2(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5490_ (.A1(_0655_),
    .A2(_0666_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5491_ (.A1(_0641_),
    .A2(_0645_),
    .A3(_0667_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5492_ (.A1(_0625_),
    .A2(_0668_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5493_ (.A1(_0622_),
    .A2(_0669_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5494_ (.A1(_0601_),
    .A2(_0670_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5495_ (.A1(_0599_),
    .A2(_0671_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5496_ (.A1(_0587_),
    .A2(_0672_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5497_ (.A1(_0587_),
    .A2(_0672_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5498_ (.A1(_0451_),
    .A2(_0673_),
    .B(_0674_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5499_ (.I(_0598_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5500_ (.A1(_0595_),
    .A2(_0596_),
    .B(_0594_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5501_ (.A1(_0588_),
    .A2(_0676_),
    .B(_0677_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5502_ (.A1(_0546_),
    .A2(_0583_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5503_ (.A1(_0600_),
    .A2(_0679_),
    .B(_0670_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5504_ (.A1(_0599_),
    .A2(_0671_),
    .B(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5505_ (.A1(_0589_),
    .A2(_0593_),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5506_ (.A1(_0606_),
    .A2(_0620_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5507_ (.A1(_0604_),
    .A2(_0621_),
    .B(_0683_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5508_ (.A1(_0590_),
    .A2(_0609_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5509_ (.A1(_0608_),
    .A2(_0610_),
    .B(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5510_ (.I(_0444_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5511_ (.A1(_0027_),
    .A2(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5512_ (.A1(_0686_),
    .A2(_0688_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5513_ (.A1(_0686_),
    .A2(_0688_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5514_ (.A1(_0689_),
    .A2(_0690_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5515_ (.A1(_0684_),
    .A2(_0691_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5516_ (.A1(_0682_),
    .A2(_0692_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5517_ (.A1(_0625_),
    .A2(_0668_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5518_ (.A1(_0622_),
    .A2(_0669_),
    .B(_0694_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5519_ (.A1(_0645_),
    .A2(_0667_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5520_ (.A1(_0645_),
    .A2(_0667_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5521_ (.A1(_0641_),
    .A2(_0696_),
    .B(_0697_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5522_ (.A1(_0637_),
    .A2(_0638_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5523_ (.A1(_0637_),
    .A2(_0638_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5524_ (.A1(_0699_),
    .A2(_0639_),
    .B(_0700_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5525_ (.A1(_3922_),
    .A2(_3772_),
    .A3(_0646_),
    .A4(_0651_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5526_ (.A1(_0652_),
    .A2(_0654_),
    .B(_0702_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5527_ (.A1(_4010_),
    .A2(_0401_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5528_ (.A1(_4015_),
    .A2(_0393_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5529_ (.A1(_0703_),
    .A2(_0704_),
    .A3(_0705_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5530_ (.A1(_0701_),
    .A2(_0706_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5531_ (.A1(_0661_),
    .A2(_0665_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5532_ (.A1(_0655_),
    .A2(_0666_),
    .B(_0708_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5533_ (.I(_0656_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5534_ (.I(_0710_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5535_ (.A1(_3973_),
    .A2(\C[2][9] ),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5536_ (.A1(_4198_),
    .A2(_0711_),
    .A3(_0712_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5537_ (.A1(_4198_),
    .A2(_0711_),
    .B1(_0712_),
    .B2(_0469_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5538_ (.A1(_0713_),
    .A2(_0714_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5539_ (.I(_0648_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5540_ (.A1(_4273_),
    .A2(_0716_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5541_ (.I(_0646_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5542_ (.A1(_4218_),
    .A2(_0718_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5543_ (.I(_0571_),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5544_ (.A1(_4169_),
    .A2(_0720_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5545_ (.A1(_0717_),
    .A2(_0719_),
    .A3(_0721_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5546_ (.A1(_0663_),
    .A2(_0715_),
    .A3(_0722_),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5547_ (.A1(_0707_),
    .A2(_0709_),
    .A3(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5548_ (.I(_0614_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5549_ (.A1(_0725_),
    .A2(_0618_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5550_ (.A1(_0611_),
    .A2(_0619_),
    .B(_0726_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5551_ (.A1(_0636_),
    .A2(_0640_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5552_ (.A1(_0636_),
    .A2(_0640_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5553_ (.A1(_0629_),
    .A2(_0728_),
    .B(_0729_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5554_ (.A1(_3842_),
    .A2(_0409_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5555_ (.A1(_3304_),
    .A2(_0319_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5556_ (.A1(_3615_),
    .A2(_0529_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5557_ (.A1(_0732_),
    .A2(_0733_),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5558_ (.A1(_0731_),
    .A2(_0734_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5559_ (.A1(_0574_),
    .A2(_0537_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5560_ (.A1(_4061_),
    .A2(_0539_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5561_ (.A1(_0512_),
    .A2(_0537_),
    .B1(_0539_),
    .B2(_4015_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5562_ (.A1(_0512_),
    .A2(_4015_),
    .A3(_0537_),
    .A4(_0533_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5563_ (.A1(_0738_),
    .A2(_0617_),
    .B(_0739_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5564_ (.A1(_0736_),
    .A2(_0737_),
    .A3(_0740_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5565_ (.A1(_0735_),
    .A2(_0741_),
    .Z(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5566_ (.A1(_0730_),
    .A2(_0742_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5567_ (.A1(_0727_),
    .A2(_0743_),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5568_ (.A1(_0698_),
    .A2(_0724_),
    .A3(_0744_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5569_ (.A1(_0695_),
    .A2(_0745_),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5570_ (.A1(_0693_),
    .A2(_0746_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5571_ (.A1(_0678_),
    .A2(_0681_),
    .A3(_0747_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5572_ (.A1(_0675_),
    .A2(_0748_),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5573_ (.I(_0320_),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5574_ (.I(_0750_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5575_ (.I(_0313_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5576_ (.I(_0751_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5577_ (.A1(_0207_),
    .A2(_0752_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5578_ (.A1(_0201_),
    .A2(_0052_),
    .A3(_0753_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5579_ (.A1(\A[2][5] ),
    .A2(_4078_),
    .B1(_3271_),
    .B2(_4077_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5580_ (.A1(_3822_),
    .A2(_0755_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5581_ (.I(_0756_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5582_ (.I(_0436_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5583_ (.A1(_0021_),
    .A2(_0757_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5584_ (.A1(_0754_),
    .A2(_0758_),
    .Z(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5585_ (.A1(_3876_),
    .A2(_0315_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5586_ (.I(_0317_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5587_ (.A1(_0206_),
    .A2(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5588_ (.A1(_0760_),
    .A2(_0762_),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5589_ (.A1(_0199_),
    .A2(_0345_),
    .B1(_0415_),
    .B2(_0386_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5590_ (.I(_0423_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5591_ (.A1(_0356_),
    .A2(_0033_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5592_ (.A1(_0489_),
    .A2(_0199_),
    .A3(_0345_),
    .A4(_0415_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5593_ (.A1(_0764_),
    .A2(_0765_),
    .B(_0766_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5594_ (.A1(_2889_),
    .A2(_0363_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5595_ (.A1(_3772_),
    .A2(_0354_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5596_ (.A1(_0768_),
    .A2(_0769_),
    .A3(_0361_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5597_ (.A1(_0767_),
    .A2(_0770_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5598_ (.A1(_0767_),
    .A2(_0770_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5599_ (.A1(_0763_),
    .A2(_0771_),
    .B(_0772_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5600_ (.I(_3964_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5601_ (.I(_0389_),
    .Z(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5602_ (.A1(_0774_),
    .A2(_0203_),
    .A3(_0378_),
    .A4(_0775_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5603_ (.A1(_2706_),
    .A2(_0493_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5604_ (.A1(_3814_),
    .A2(_0383_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5605_ (.A1(_0777_),
    .A2(_0778_),
    .A3(_0394_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5606_ (.A1(_0776_),
    .A2(_0779_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5607_ (.A1(_0309_),
    .A2(_0316_),
    .A3(_0321_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5608_ (.A1(_0366_),
    .A2(_0370_),
    .A3(_0781_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5609_ (.A1(_0780_),
    .A2(_0782_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5610_ (.A1(_0780_),
    .A2(_0782_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5611_ (.A1(_0773_),
    .A2(_0783_),
    .B(_0784_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5612_ (.A1(_0022_),
    .A2(_0436_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5613_ (.A1(_0329_),
    .A2(_0786_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5614_ (.A1(_0785_),
    .A2(_0787_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5615_ (.A1(_0759_),
    .A2(_0788_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5616_ (.A1(_0773_),
    .A2(_0783_),
    .Z(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5617_ (.A1(_0776_),
    .A2(_0779_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5618_ (.A1(_0465_),
    .A2(_0470_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5619_ (.A1(_3973_),
    .A2(\C[2][2] ),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5620_ (.A1(_0342_),
    .A2(_0498_),
    .A3(_0793_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5621_ (.I(_0476_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5622_ (.A1(_0795_),
    .A2(_0458_),
    .B1(_0466_),
    .B2(_2717_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5623_ (.A1(_0794_),
    .A2(_0796_),
    .B(_0463_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5624_ (.A1(_0792_),
    .A2(_0797_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5625_ (.A1(_4198_),
    .A2(_0462_),
    .A3(_0793_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5626_ (.I(_3845_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5627_ (.A1(_0800_),
    .A2(_0458_),
    .A3(_0466_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5628_ (.A1(_0801_),
    .A2(_0796_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5629_ (.A1(_0792_),
    .A2(_0799_),
    .A3(_0802_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5630_ (.A1(_0791_),
    .A2(_0798_),
    .B(_0803_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5631_ (.A1(_0471_),
    .A2(_0483_),
    .A3(_0455_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5632_ (.A1(_0804_),
    .A2(_0805_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5633_ (.A1(_0804_),
    .A2(_0805_),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5634_ (.A1(_0790_),
    .A2(_0806_),
    .B(_0807_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5635_ (.A1(_0486_),
    .A2(_0521_),
    .A3(_0454_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5636_ (.A1(_0808_),
    .A2(_0809_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5637_ (.A1(_0808_),
    .A2(_0809_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5638_ (.A1(_0789_),
    .A2(_0810_),
    .B(_0811_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5639_ (.A1(_0452_),
    .A2(_0585_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5640_ (.A1(_0812_),
    .A2(_0813_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5641_ (.A1(_0785_),
    .A2(_0787_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5642_ (.A1(_0759_),
    .A2(_0788_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5643_ (.A1(_0815_),
    .A2(_0816_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5644_ (.A1(_0453_),
    .A2(_0585_),
    .A3(_0812_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5645_ (.A1(_0817_),
    .A2(_0818_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5646_ (.A1(_0587_),
    .A2(_0672_),
    .A3(_0451_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5647_ (.A1(_0814_),
    .A2(_0819_),
    .B(_0820_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5648_ (.I(_0345_),
    .Z(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5649_ (.A1(_0347_),
    .A2(_0351_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5650_ (.I(_0822_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5651_ (.A1(_3871_),
    .A2(_0050_),
    .B1(_0823_),
    .B2(_4275_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5652_ (.A1(_0489_),
    .A2(_0033_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5653_ (.A1(_4275_),
    .A2(_3871_),
    .A3(_0414_),
    .A4(_0823_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5654_ (.A1(_0824_),
    .A2(_0825_),
    .B(_0826_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5655_ (.A1(_3875_),
    .A2(_0364_),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5656_ (.A1(_0386_),
    .A2(_0533_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5657_ (.A1(_0828_),
    .A2(_0829_),
    .A3(_0765_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5658_ (.A1(_0827_),
    .A2(_0830_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5659_ (.A1(_0827_),
    .A2(_0830_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5660_ (.A1(_0753_),
    .A2(_0831_),
    .B(_0832_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5661_ (.A1(_0763_),
    .A2(_0771_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5662_ (.A1(_0833_),
    .A2(_0834_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5663_ (.A1(_0754_),
    .A2(_0758_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5664_ (.A1(_0833_),
    .A2(_0834_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5665_ (.I(_0377_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5666_ (.A1(_0203_),
    .A2(_0838_),
    .B1(_0775_),
    .B2(_0774_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5667_ (.I(_0839_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5668_ (.A1(_0776_),
    .A2(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5669_ (.A1(_3973_),
    .A2(\C[2][1] ),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5670_ (.A1(_0199_),
    .A2(_0498_),
    .A3(_0842_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5671_ (.A1(_0342_),
    .A2(_0498_),
    .B1(_0793_),
    .B2(_0795_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5672_ (.A1(_0843_),
    .A2(_0844_),
    .B(_0794_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5673_ (.A1(_0802_),
    .A2(_0845_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5674_ (.A1(_0200_),
    .A2(_0467_),
    .A3(_0842_),
    .Z(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5675_ (.A1(_0799_),
    .A2(_0844_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5676_ (.A1(_0802_),
    .A2(_0847_),
    .A3(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5677_ (.A1(_0841_),
    .A2(_0846_),
    .B(_0849_),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5678_ (.A1(_0791_),
    .A2(_0798_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5679_ (.A1(_0850_),
    .A2(_0851_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5680_ (.A1(_0850_),
    .A2(_0851_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5681_ (.A1(_0837_),
    .A2(_0852_),
    .B(_0853_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5682_ (.A1(_0790_),
    .A2(_0806_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5683_ (.A1(_0854_),
    .A2(_0855_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5684_ (.A1(_0835_),
    .A2(_0836_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5685_ (.I(_0857_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5686_ (.A1(_0854_),
    .A2(_0855_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5687_ (.A1(_0858_),
    .A2(_0859_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5688_ (.A1(_0789_),
    .A2(_0810_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5689_ (.A1(_0856_),
    .A2(_0860_),
    .A3(_0861_),
    .ZN(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5690_ (.A1(_0856_),
    .A2(_0860_),
    .B(_0861_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5691_ (.A1(_0835_),
    .A2(_0836_),
    .A3(_0862_),
    .B(_0863_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5692_ (.A1(_0817_),
    .A2(_0818_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5693_ (.A1(_0864_),
    .A2(_0865_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5694_ (.A1(_0857_),
    .A2(_0859_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5695_ (.A1(_0020_),
    .A2(_0757_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5696_ (.I(_0868_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5697_ (.A1(_0753_),
    .A2(_0831_),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5698_ (.A1(\C[2][0] ),
    .A2(_3870_),
    .A3(_4239_),
    .A4(_0462_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5699_ (.I(_0871_),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5700_ (.A1(_3876_),
    .A2(_0462_),
    .B1(_0842_),
    .B2(_0795_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5701_ (.A1(_0847_),
    .A2(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5702_ (.A1(_0848_),
    .A2(_0874_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5703_ (.A1(_0200_),
    .A2(_0838_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5704_ (.A1(_0871_),
    .A2(_0873_),
    .B(_0843_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5705_ (.A1(_0848_),
    .A2(_0877_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5706_ (.A1(_0872_),
    .A2(_0875_),
    .B1(_0876_),
    .B2(_0878_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5707_ (.A1(_0841_),
    .A2(_0846_),
    .Z(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5708_ (.A1(_0879_),
    .A2(_0880_),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5709_ (.A1(_0879_),
    .A2(_0880_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5710_ (.A1(_0870_),
    .A2(_0881_),
    .B(_0882_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5711_ (.A1(_0850_),
    .A2(_0851_),
    .A3(_0837_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5712_ (.A1(_0883_),
    .A2(_0884_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5713_ (.A1(_0883_),
    .A2(_0884_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5714_ (.A1(_0869_),
    .A2(_0885_),
    .B(_0886_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5715_ (.A1(_0867_),
    .A2(_0887_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5716_ (.A1(_0835_),
    .A2(_0836_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5717_ (.A1(_0858_),
    .A2(_0859_),
    .B(_0856_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5718_ (.A1(_0889_),
    .A2(_0890_),
    .A3(_0861_),
    .Z(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5719_ (.A1(_0888_),
    .A2(_0891_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5720_ (.I(_0892_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5721_ (.A1(_0336_),
    .A2(_0334_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5722_ (.I(_0894_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5723_ (.A1(_4073_),
    .A2(_0032_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5724_ (.I(_0343_),
    .Z(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5725_ (.I(_0896_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5726_ (.A1(_0206_),
    .A2(_0897_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5727_ (.I(_0823_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5728_ (.A1(_0774_),
    .A2(_0899_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5729_ (.A1(_0898_),
    .A2(_0900_),
    .A3(_0825_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5730_ (.I(_0901_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5731_ (.I(_0493_),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5732_ (.A1(_0847_),
    .A2(_0871_),
    .A3(_0873_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5733_ (.A1(_0847_),
    .A2(_0873_),
    .B(_0872_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5734_ (.A1(_3882_),
    .A2(_0903_),
    .A3(_0904_),
    .A4(_0905_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5735_ (.A1(_0848_),
    .A2(_0876_),
    .A3(_0877_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5736_ (.A1(_0906_),
    .A2(_0907_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5737_ (.A1(_0906_),
    .A2(_0907_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5738_ (.A1(_0902_),
    .A2(_0908_),
    .B(_0909_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5739_ (.A1(_0879_),
    .A2(_0880_),
    .A3(_0870_),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5740_ (.A1(_0910_),
    .A2(_0911_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5741_ (.A1(_0910_),
    .A2(_0911_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5742_ (.A1(_0895_),
    .A2(_0912_),
    .B(_0913_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5743_ (.A1(_0883_),
    .A2(_0884_),
    .A3(_0869_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5744_ (.A1(_0914_),
    .A2(_0915_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5745_ (.A1(_0867_),
    .A2(_0887_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5746_ (.A1(_0888_),
    .A2(_0916_),
    .A3(_0917_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _5747_ (.A1(_0910_),
    .A2(_0911_),
    .A3(_0895_),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5748_ (.I(_0334_),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5749_ (.A1(_0336_),
    .A2(_3790_),
    .A3(_0920_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5750_ (.I(_0774_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5751_ (.I(_0358_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5752_ (.I(_0359_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5753_ (.A1(_0922_),
    .A2(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5754_ (.I(_0924_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5755_ (.I(_0903_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5756_ (.A1(_0024_),
    .A2(_0049_),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5757_ (.A1(_0872_),
    .A2(_0874_),
    .A3(_0926_),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5758_ (.A1(_0016_),
    .A2(_0925_),
    .A3(_0927_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5759_ (.A1(_0906_),
    .A2(_0907_),
    .A3(_0902_),
    .Z(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5760_ (.A1(_0928_),
    .A2(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5761_ (.A1(_0928_),
    .A2(_0929_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5762_ (.A1(_0921_),
    .A2(_0930_),
    .B(_0931_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5763_ (.A1(_0914_),
    .A2(_0915_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5764_ (.A1(_0916_),
    .A2(_0919_),
    .A3(_0932_),
    .A4(_0933_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5765_ (.A1(_0919_),
    .A2(_0932_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5766_ (.A1(_0919_),
    .A2(_0932_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5767_ (.I(_0336_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5768_ (.A1(_0016_),
    .A2(_0925_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5769_ (.A1(_0927_),
    .A2(_0938_),
    .Z(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5770_ (.A1(_0937_),
    .A2(_0181_),
    .A3(_0920_),
    .A4(_0939_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5771_ (.A1(_0928_),
    .A2(_0929_),
    .A3(_0921_),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5772_ (.A1(_0940_),
    .A2(_0941_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5773_ (.A1(_0937_),
    .A2(_0181_),
    .A3(_0920_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5774_ (.A1(_0939_),
    .A2(_0943_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5775_ (.I(_0467_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5776_ (.I(_0945_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5777_ (.A1(_0024_),
    .A2(_0048_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5778_ (.I(_0186_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5779_ (.A1(\C[2][0] ),
    .A2(_0947_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5780_ (.A1(_0946_),
    .A2(_0948_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5781_ (.A1(_0872_),
    .A2(_0949_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5782_ (.A1(_0016_),
    .A2(_0757_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5783_ (.A1(_0950_),
    .A2(_0951_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5784_ (.A1(_0944_),
    .A2(_0952_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5785_ (.A1(_0941_),
    .A2(_0953_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5786_ (.A1(_0919_),
    .A2(_0932_),
    .A3(_0942_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5787_ (.A1(_0935_),
    .A2(_0936_),
    .A3(_0942_),
    .B1(_0954_),
    .B2(_0955_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5788_ (.A1(_0914_),
    .A2(_0915_),
    .A3(_0935_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5789_ (.A1(_0956_),
    .A2(_0957_),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5790_ (.A1(_0867_),
    .A2(_0887_),
    .A3(_0916_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5791_ (.A1(_0934_),
    .A2(_0958_),
    .B(_0959_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5792_ (.A1(_0888_),
    .A2(_0891_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5793_ (.A1(_0918_),
    .A2(_0960_),
    .B(_0961_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5794_ (.A1(_0864_),
    .A2(_0865_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5795_ (.A1(_0893_),
    .A2(_0962_),
    .B(_0963_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5796_ (.A1(_0866_),
    .A2(_0964_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5797_ (.A1(_0814_),
    .A2(_0819_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5798_ (.A1(_0966_),
    .A2(_0820_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5799_ (.A1(_0965_),
    .A2(_0967_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5800_ (.A1(_0821_),
    .A2(_0968_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5801_ (.A1(_0749_),
    .A2(_0969_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5802_ (.I(_0970_),
    .Z(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5803_ (.A1(_4105_),
    .A2(_4192_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5804_ (.A1(_3911_),
    .A2(_4193_),
    .B(_0971_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5805_ (.I(_0220_),
    .Z(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5806_ (.A1(_4107_),
    .A2(_0057_),
    .A3(_4115_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5807_ (.I(_4107_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5808_ (.A1(_0031_),
    .A2(_0057_),
    .B(_4115_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _5809_ (.A1(_4111_),
    .A2(_0973_),
    .A3(_0974_),
    .B1(_4119_),
    .B2(_4109_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5810_ (.A1(_4122_),
    .A2(_4190_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5811_ (.A1(_4120_),
    .A2(_4191_),
    .B(_0976_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5812_ (.A1(_4127_),
    .A2(_4144_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5813_ (.A1(_4124_),
    .A2(_4145_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5814_ (.I(_3026_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5815_ (.I(_3315_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5816_ (.A1(_0980_),
    .A2(_0981_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5817_ (.A1(_4128_),
    .A2(_4131_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5818_ (.A1(_4028_),
    .A2(_0982_),
    .B1(_0983_),
    .B2(_4129_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5819_ (.A1(_0978_),
    .A2(_0979_),
    .B(_0984_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5820_ (.A1(_0978_),
    .A2(_0979_),
    .A3(_0984_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5821_ (.A1(_0985_),
    .A2(_0986_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5822_ (.A1(_0973_),
    .A2(_0987_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5823_ (.A1(_4165_),
    .A2(_4188_),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5824_ (.A1(_4165_),
    .A2(_4188_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5825_ (.A1(_4149_),
    .A2(_4189_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5826_ (.I(_4146_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5827_ (.A1(_4149_),
    .A2(_0989_),
    .A3(_0990_),
    .B1(_0991_),
    .B2(_0992_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5828_ (.A1(_4139_),
    .A2(_4142_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5829_ (.A1(_4132_),
    .A2(_4143_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5830_ (.A1(_0994_),
    .A2(_0995_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5831_ (.A1(_4156_),
    .A2(_4163_),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5832_ (.A1(_4153_),
    .A2(_4164_),
    .B(_0997_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5833_ (.A1(_2460_),
    .A2(_3897_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5834_ (.A1(_3849_),
    .A2(_3615_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5835_ (.A1(_0982_),
    .A2(_0999_),
    .A3(_1000_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5836_ (.A1(_0310_),
    .A2(_4137_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5837_ (.A1(_4136_),
    .A2(_4141_),
    .Z(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5838_ (.A1(_3868_),
    .A2(_1002_),
    .B1(_1003_),
    .B2(_4140_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5839_ (.A1(_0397_),
    .A2(_3863_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5840_ (.A1(_0800_),
    .A2(_3873_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5841_ (.A1(_1002_),
    .A2(_1005_),
    .A3(_1006_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5842_ (.A1(_1004_),
    .A2(_1007_),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5843_ (.A1(_1001_),
    .A2(_1008_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5844_ (.A1(_0998_),
    .A2(_1009_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5845_ (.A1(_0996_),
    .A2(_1010_),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5846_ (.A1(_4167_),
    .A2(_4187_),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5847_ (.A1(_4165_),
    .A2(_4188_),
    .B(_1012_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5848_ (.A1(_4181_),
    .A2(_4183_),
    .A3(_4185_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5849_ (.A1(_4181_),
    .A2(_4183_),
    .B(_4185_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5850_ (.A1(_4178_),
    .A2(_1014_),
    .A3(_1015_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5851_ (.A1(_4175_),
    .A2(_4186_),
    .B(_1016_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5852_ (.I(_3934_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5853_ (.A1(_3761_),
    .A2(_4168_),
    .A3(_1018_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5854_ (.I(_0755_),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5855_ (.A1(_4001_),
    .A2(_3948_),
    .A3(_1020_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5856_ (.A1(_1019_),
    .A2(_1021_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5857_ (.A1(_0043_),
    .A2(_0541_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5858_ (.A1(_1022_),
    .A2(_1023_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5859_ (.A1(_3822_),
    .A2(_3824_),
    .A3(_4179_),
    .A4(_4180_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5860_ (.A1(_4183_),
    .A2(_4185_),
    .B(_1025_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5861_ (.A1(_0513_),
    .A2(\C[3][9] ),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _5862_ (.A1(_3777_),
    .A2(_3789_),
    .A3(_4182_),
    .A4(_1027_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _5863_ (.A1(_3777_),
    .A2(_3789_),
    .A3(_4182_),
    .B1(_1027_),
    .B2(_3926_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5864_ (.A1(_1028_),
    .A2(_1029_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5865_ (.A1(_4045_),
    .A2(_4067_),
    .A3(_4096_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5866_ (.A1(_1026_),
    .A2(_1030_),
    .A3(_1031_),
    .Z(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5867_ (.A1(_1024_),
    .A2(_1032_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5868_ (.A1(_1017_),
    .A2(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5869_ (.A1(_4069_),
    .A2(_0020_),
    .A3(_4068_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5870_ (.A1(_4171_),
    .A2(_4174_),
    .B(_1035_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5871_ (.I(_4062_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5872_ (.I(_1037_),
    .Z(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5873_ (.A1(_4160_),
    .A2(_4162_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5874_ (.A1(_0042_),
    .A2(_1038_),
    .A3(_1039_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5875_ (.A1(_1036_),
    .A2(_1040_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5876_ (.A1(_1034_),
    .A2(_1041_),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5877_ (.A1(_1013_),
    .A2(_1042_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5878_ (.A1(_1011_),
    .A2(_1043_),
    .Z(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5879_ (.A1(_0988_),
    .A2(_0993_),
    .A3(_1044_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5880_ (.A1(_0975_),
    .A2(_0977_),
    .A3(_1045_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5881_ (.A1(_0972_),
    .A2(_1046_),
    .Z(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5882_ (.A1(_4194_),
    .A2(_4260_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5883_ (.A1(_4261_),
    .A2(_0301_),
    .B(_1048_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5884_ (.A1(_1047_),
    .A2(_1049_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5885_ (.I(_1050_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5886_ (.A1(_0589_),
    .A2(_0593_),
    .A3(_0692_),
    .B1(_0691_),
    .B2(_0684_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5887_ (.A1(_0695_),
    .A2(_0745_),
    .Z(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5888_ (.A1(_0693_),
    .A2(_0746_),
    .B(_1052_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5889_ (.A1(_0730_),
    .A2(_0742_),
    .Z(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5890_ (.A1(_0727_),
    .A2(_0743_),
    .B(_1054_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5891_ (.A1(_3625_),
    .A2(_0750_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5892_ (.I(_1056_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5893_ (.A1(_0609_),
    .A2(_1057_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5894_ (.A1(_0731_),
    .A2(_0734_),
    .B(_1058_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5895_ (.A1(_0028_),
    .A2(_0445_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5896_ (.A1(_1059_),
    .A2(_1060_),
    .Z(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5897_ (.A1(_1059_),
    .A2(_1060_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5898_ (.A1(_1061_),
    .A2(_1062_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5899_ (.A1(_1055_),
    .A2(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5900_ (.A1(_0689_),
    .A2(_1064_),
    .Z(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5901_ (.A1(_0698_),
    .A2(_0724_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5902_ (.I(_0744_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5903_ (.A1(_0698_),
    .A2(_0724_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5904_ (.A1(_1066_),
    .A2(_1067_),
    .B(_1068_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5905_ (.A1(_0736_),
    .A2(_0737_),
    .Z(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5906_ (.A1(_0736_),
    .A2(_0737_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5907_ (.A1(_1070_),
    .A2(_1071_),
    .A3(_0740_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5908_ (.A1(_0735_),
    .A2(_0741_),
    .B(_1072_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5909_ (.A1(_0704_),
    .A2(_0705_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5910_ (.A1(_0704_),
    .A2(_0705_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5911_ (.A1(_0703_),
    .A2(_1074_),
    .A3(_1075_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5912_ (.A1(_0701_),
    .A2(_0706_),
    .B(_1076_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5913_ (.A1(_4026_),
    .A2(_0409_),
    .Z(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5914_ (.A1(_3897_),
    .A2(_0051_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5915_ (.A1(_1056_),
    .A2(_1078_),
    .A3(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5916_ (.A1(_1070_),
    .A2(_1080_),
    .Z(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5917_ (.A1(_1077_),
    .A2(_1081_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5918_ (.A1(_1073_),
    .A2(_1082_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5919_ (.A1(_0709_),
    .A2(_0723_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5920_ (.A1(_0709_),
    .A2(_0723_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5921_ (.A1(_0707_),
    .A2(_1084_),
    .B(_1085_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5922_ (.A1(_4218_),
    .A2(_0647_),
    .B1(_0649_),
    .B2(_3773_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5923_ (.A1(_4218_),
    .A2(_4273_),
    .A3(_0647_),
    .A4(_0649_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5924_ (.A1(_1087_),
    .A2(_0721_),
    .B(_1088_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5925_ (.A1(_0541_),
    .A2(_0488_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5926_ (.A1(_1037_),
    .A2(_0403_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5927_ (.A1(_1089_),
    .A2(_1090_),
    .A3(_1091_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5928_ (.A1(_1074_),
    .A2(_1092_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5929_ (.I(_0657_),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5930_ (.A1(_3876_),
    .A2(_1094_),
    .A3(_0662_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5931_ (.A1(_0713_),
    .A2(_0714_),
    .B(_1095_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5932_ (.A1(_1095_),
    .A2(_0713_),
    .A3(_0714_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5933_ (.A1(_1096_),
    .A2(_0722_),
    .B(_1097_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5934_ (.I(_0657_),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5935_ (.A1(_0342_),
    .A2(_1099_),
    .A3(_0712_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5936_ (.A1(_3983_),
    .A2(\C[2][10] ),
    .Z(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5937_ (.A1(_0800_),
    .A2(_0710_),
    .A3(_1101_),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5938_ (.A1(_0800_),
    .A2(_0710_),
    .B1(_1101_),
    .B2(_3976_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5939_ (.A1(_1102_),
    .A2(_1103_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5940_ (.A1(_4072_),
    .A2(_0649_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5941_ (.A1(_3805_),
    .A2(_0646_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5942_ (.A1(_0422_),
    .A2(_0720_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5943_ (.A1(_1105_),
    .A2(_1106_),
    .A3(_1107_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5944_ (.A1(_1100_),
    .A2(_1104_),
    .A3(_1108_),
    .Z(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5945_ (.A1(_1098_),
    .A2(_1109_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5946_ (.A1(_1093_),
    .A2(_1110_),
    .Z(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5947_ (.A1(_1086_),
    .A2(_1111_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5948_ (.A1(_1083_),
    .A2(_1112_),
    .Z(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5949_ (.A1(_1065_),
    .A2(_1069_),
    .A3(_1113_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5950_ (.A1(_1053_),
    .A2(_1114_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5951_ (.A1(_1051_),
    .A2(_1115_),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5952_ (.A1(_0681_),
    .A2(_0747_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5953_ (.A1(_0681_),
    .A2(_0747_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5954_ (.A1(_0678_),
    .A2(_1117_),
    .B(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5955_ (.A1(_1116_),
    .A2(_1119_),
    .Z(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5956_ (.A1(_0866_),
    .A2(_0964_),
    .B(_0967_),
    .C(_0749_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5957_ (.A1(_0675_),
    .A2(_0748_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5958_ (.A1(_0675_),
    .A2(_0748_),
    .B(_0821_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5959_ (.A1(_1122_),
    .A2(_1123_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5960_ (.A1(_1121_),
    .A2(_1124_),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5961_ (.A1(_1120_),
    .A2(_1125_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5962_ (.I(_1126_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5963_ (.A1(_0973_),
    .A2(_0987_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5964_ (.A1(_0985_),
    .A2(_1127_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5965_ (.A1(_0993_),
    .A2(_1044_),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5966_ (.A1(_0993_),
    .A2(_1044_),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5967_ (.A1(_0988_),
    .A2(_1129_),
    .B(_1130_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5968_ (.A1(_0998_),
    .A2(_1009_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5969_ (.A1(_0994_),
    .A2(_0995_),
    .B(_1010_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5970_ (.A1(_1132_),
    .A2(_1133_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5971_ (.I(_0980_),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5972_ (.A1(_0060_),
    .A2(_0030_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5973_ (.A1(_0982_),
    .A2(_1000_),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5974_ (.A1(_4131_),
    .A2(_1135_),
    .B1(_1136_),
    .B2(_0999_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5975_ (.A1(_1134_),
    .A2(_1137_),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5976_ (.A1(_1012_),
    .A2(_0989_),
    .B(_1042_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5977_ (.A1(_1011_),
    .A2(_1043_),
    .B(_1139_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5978_ (.A1(_1004_),
    .A2(_1007_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5979_ (.A1(_1001_),
    .A2(_1008_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5980_ (.A1(_1141_),
    .A2(_1142_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5981_ (.A1(_4215_),
    .A2(_4159_),
    .A3(_1036_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5982_ (.A1(_1039_),
    .A2(_1144_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5983_ (.A1(_3844_),
    .A2(_0574_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5984_ (.A1(_1000_),
    .A2(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5985_ (.A1(_4195_),
    .A2(_3897_),
    .B1(_3625_),
    .B2(_4202_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5986_ (.A1(_1147_),
    .A2(_1148_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5987_ (.A1(_2685_),
    .A2(_4135_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5988_ (.A1(_2695_),
    .A2(_3872_),
    .B1(_4137_),
    .B2(_4031_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5989_ (.A1(_4141_),
    .A2(_1150_),
    .B1(_1151_),
    .B2(_1005_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5990_ (.A1(_3862_),
    .A2(_3293_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5991_ (.A1(_0397_),
    .A2(_3867_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5992_ (.A1(_1150_),
    .A2(_1153_),
    .A3(_1154_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5993_ (.A1(_1152_),
    .A2(_1155_),
    .Z(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5994_ (.A1(_1149_),
    .A2(_1156_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5995_ (.I(_1157_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5996_ (.A1(_1145_),
    .A2(_1158_),
    .Z(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5997_ (.A1(_1143_),
    .A2(_1159_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5998_ (.A1(_1017_),
    .A2(_1033_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5999_ (.A1(_1034_),
    .A2(_1041_),
    .B(_1161_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6000_ (.A1(_3916_),
    .A2(_3760_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6001_ (.I(_1163_),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6002_ (.A1(_1164_),
    .A2(_1020_),
    .A3(_1019_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6003_ (.A1(_1022_),
    .A2(_1023_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6004_ (.A1(_1165_),
    .A2(_1166_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6005_ (.A1(_1028_),
    .A2(_1029_),
    .A3(_1031_),
    .Z(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6006_ (.A1(_1028_),
    .A2(_1029_),
    .B(_1031_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6007_ (.A1(_1026_),
    .A2(_1168_),
    .A3(_1169_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6008_ (.A1(_1024_),
    .A2(_1032_),
    .B(_1170_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6009_ (.A1(_4172_),
    .A2(_4062_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6010_ (.A1(_0021_),
    .A2(_3998_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6011_ (.A1(_1164_),
    .A2(_0337_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6012_ (.A1(_1172_),
    .A2(_1173_),
    .A3(_1174_),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6013_ (.A1(_3993_),
    .A2(_3790_),
    .A3(_4093_),
    .A4(_1027_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6014_ (.A1(_1029_),
    .A2(_1031_),
    .B(_1176_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6015_ (.I(_3890_),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6016_ (.A1(_1178_),
    .A2(\C[3][10] ),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _6017_ (.A1(_4045_),
    .A2(_4067_),
    .A3(_4179_),
    .A4(_1179_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6018_ (.I(_3925_),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _6019_ (.A1(_4045_),
    .A2(_4067_),
    .A3(_4093_),
    .B1(_1179_),
    .B2(_1181_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6020_ (.A1(_1180_),
    .A2(_1182_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6021_ (.I(_3992_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6022_ (.A1(_1184_),
    .A2(_4080_),
    .A3(_4096_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6023_ (.A1(_1177_),
    .A2(_1183_),
    .A3(_1185_),
    .Z(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6024_ (.A1(_1175_),
    .A2(_1186_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6025_ (.A1(_1171_),
    .A2(_1187_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6026_ (.A1(_1167_),
    .A2(_1188_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6027_ (.A1(_1160_),
    .A2(_1162_),
    .A3(_1189_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6028_ (.A1(_1140_),
    .A2(_1190_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6029_ (.A1(_1138_),
    .A2(_1191_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6030_ (.A1(_1131_),
    .A2(_1192_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6031_ (.A1(_1128_),
    .A2(_1193_),
    .Z(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6032_ (.A1(_0977_),
    .A2(_1045_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6033_ (.A1(_0977_),
    .A2(_1045_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6034_ (.A1(_0975_),
    .A2(_1195_),
    .B(_1196_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6035_ (.A1(_1194_),
    .A2(_1197_),
    .Z(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6036_ (.A1(_4261_),
    .A2(_0178_),
    .A3(_0300_),
    .A4(_1047_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6037_ (.A1(_0972_),
    .A2(_1046_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6038_ (.A1(_0972_),
    .A2(_1046_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6039_ (.A1(_1048_),
    .A2(_1200_),
    .B(_1201_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6040_ (.A1(_1199_),
    .A2(_1202_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6041_ (.A1(_1198_),
    .A2(_1203_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6042_ (.I(_1204_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6043_ (.A1(_1053_),
    .A2(_1114_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6044_ (.A1(_1051_),
    .A2(_1115_),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6045_ (.A1(_1055_),
    .A2(_1063_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6046_ (.A1(_0689_),
    .A2(_1064_),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6047_ (.A1(_1207_),
    .A2(_1208_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6048_ (.I(_1209_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6049_ (.A1(_1069_),
    .A2(_1113_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6050_ (.A1(_1069_),
    .A2(_1113_),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6051_ (.A1(_1065_),
    .A2(_1211_),
    .B(_1212_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6052_ (.A1(_1077_),
    .A2(_1081_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6053_ (.A1(_1073_),
    .A2(_1082_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6054_ (.A1(_1214_),
    .A2(_1215_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6055_ (.A1(_1057_),
    .A2(_1079_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6056_ (.A1(_1057_),
    .A2(_1079_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6057_ (.A1(_1078_),
    .A2(_1217_),
    .B(_1218_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6058_ (.A1(_0029_),
    .A2(_0687_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6059_ (.A1(_1219_),
    .A2(_1220_),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6060_ (.A1(_1219_),
    .A2(_1220_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6061_ (.A1(_1221_),
    .A2(_1222_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6062_ (.A1(_1216_),
    .A2(_1223_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6063_ (.A1(_1061_),
    .A2(_1224_),
    .Z(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6064_ (.A1(_1086_),
    .A2(_1111_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6065_ (.A1(_1083_),
    .A2(_1112_),
    .B(_1226_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6066_ (.A1(_1070_),
    .A2(_1080_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6067_ (.I(_1089_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6068_ (.A1(_1090_),
    .A2(_1091_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6069_ (.A1(_1090_),
    .A2(_1091_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6070_ (.A1(_1229_),
    .A2(_1230_),
    .A3(_1231_),
    .B1(_1092_),
    .B2(_1074_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6071_ (.A1(_3898_),
    .A2(_0607_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6072_ (.A1(_1057_),
    .A2(_1233_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6073_ (.I(_0607_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6074_ (.A1(_3905_),
    .A2(_0053_),
    .B1(_0052_),
    .B2(_3899_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6075_ (.A1(_1234_),
    .A2(_1235_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6076_ (.A1(_1232_),
    .A2(_1236_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6077_ (.A1(_1228_),
    .A2(_1237_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6078_ (.I(_1238_),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6079_ (.A1(_1098_),
    .A2(_1109_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6080_ (.A1(_1093_),
    .A2(_1110_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6081_ (.A1(_1240_),
    .A2(_1241_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6082_ (.A1(_1102_),
    .A2(_1103_),
    .B(_1100_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6083_ (.A1(_1100_),
    .A2(_1102_),
    .A3(_1103_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6084_ (.A1(_1243_),
    .A2(_1108_),
    .B(_1244_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6085_ (.A1(_0374_),
    .A2(_1099_),
    .A3(_1101_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6086_ (.I(_0456_),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6087_ (.A1(_1247_),
    .A2(\C[2][11] ),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6088_ (.A1(_3842_),
    .A2(_0710_),
    .A3(_1248_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6089_ (.A1(_0419_),
    .A2(_0658_),
    .B1(_1248_),
    .B2(_0468_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6090_ (.A1(_1249_),
    .A2(_1250_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6091_ (.I(_0508_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6092_ (.I(_1252_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6093_ (.A1(_0541_),
    .A2(_0037_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6094_ (.A1(_4168_),
    .A2(_0651_),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6095_ (.A1(_3831_),
    .A2(_0569_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6096_ (.A1(_1254_),
    .A2(_1255_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6097_ (.A1(_1253_),
    .A2(_1256_),
    .Z(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6098_ (.A1(_1246_),
    .A2(_1251_),
    .A3(_1257_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6099_ (.A1(_1245_),
    .A2(_1258_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6100_ (.A1(_1105_),
    .A2(_1106_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6101_ (.A1(_1105_),
    .A2(_1106_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6102_ (.A1(_1260_),
    .A2(_1107_),
    .B(_1261_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6103_ (.A1(_1038_),
    .A2(_0036_),
    .Z(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6104_ (.A1(_0705_),
    .A2(_1263_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6105_ (.A1(_1262_),
    .A2(_1264_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6106_ (.A1(_1259_),
    .A2(_1265_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6107_ (.A1(_1242_),
    .A2(_1266_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6108_ (.A1(_1239_),
    .A2(_1267_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6109_ (.A1(_1227_),
    .A2(_1268_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6110_ (.A1(_1225_),
    .A2(_1269_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6111_ (.A1(_1210_),
    .A2(_1213_),
    .A3(_1270_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6112_ (.A1(_1205_),
    .A2(_1206_),
    .B(_1271_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6113_ (.A1(_1205_),
    .A2(_1206_),
    .A3(_1271_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6114_ (.A1(_1272_),
    .A2(_1273_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6115_ (.A1(_1116_),
    .A2(_1119_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6116_ (.A1(_1120_),
    .A2(_1125_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6117_ (.A1(_1275_),
    .A2(_1276_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6118_ (.A1(_1274_),
    .A2(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6119_ (.I(_1278_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6120_ (.A1(_1131_),
    .A2(_1192_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6121_ (.A1(_1131_),
    .A2(_1192_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6122_ (.A1(_1128_),
    .A2(_1279_),
    .B(_1280_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6123_ (.A1(_1132_),
    .A2(_1133_),
    .B(_1137_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6124_ (.A1(_1140_),
    .A2(_1190_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6125_ (.A1(_1138_),
    .A2(_1191_),
    .B(_1283_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6126_ (.A1(_1145_),
    .A2(_1158_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6127_ (.A1(_1143_),
    .A2(_1159_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6128_ (.A1(_1285_),
    .A2(_1286_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6129_ (.A1(_1147_),
    .A2(_1287_),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6130_ (.A1(_1162_),
    .A2(_1189_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6131_ (.A1(_1162_),
    .A2(_1189_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6132_ (.A1(_1160_),
    .A2(_1289_),
    .B(_1290_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6133_ (.A1(_1152_),
    .A2(_1155_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6134_ (.A1(_1149_),
    .A2(_1156_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6135_ (.A1(_1292_),
    .A2(_1293_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6136_ (.I(_4137_),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6137_ (.A1(_0419_),
    .A2(_1295_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6138_ (.A1(_1150_),
    .A2(_1154_),
    .Z(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6139_ (.A1(_1006_),
    .A2(_1296_),
    .B1(_1297_),
    .B2(_1153_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6140_ (.A1(_3883_),
    .A2(_3636_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6141_ (.A1(_3874_),
    .A2(_0981_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6142_ (.A1(_1296_),
    .A2(_1300_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6143_ (.A1(_1299_),
    .A2(_1301_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6144_ (.A1(_1298_),
    .A2(_1302_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6145_ (.A1(_1146_),
    .A2(_1303_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6146_ (.A1(_1294_),
    .A2(_1304_),
    .Z(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6147_ (.A1(_1171_),
    .A2(_1187_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6148_ (.A1(_1167_),
    .A2(_1188_),
    .B(_1306_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6149_ (.A1(_0021_),
    .A2(_3999_),
    .B(_1174_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6150_ (.A1(_4158_),
    .A2(_4003_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6151_ (.I(_1309_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6152_ (.A1(_4173_),
    .A2(_0045_),
    .A3(_1174_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6153_ (.A1(_1172_),
    .A2(_1308_),
    .B(_1310_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6154_ (.A1(_1180_),
    .A2(_1182_),
    .A3(_1185_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6155_ (.A1(_1180_),
    .A2(_1182_),
    .B(_1185_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6156_ (.A1(_1177_),
    .A2(_1312_),
    .A3(_1313_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6157_ (.A1(_1175_),
    .A2(_1186_),
    .B(_1314_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6158_ (.A1(_0045_),
    .A2(_4161_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6159_ (.I(_1164_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6160_ (.A1(_0044_),
    .A2(_4062_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6161_ (.A1(_1316_),
    .A2(_1317_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6162_ (.I(_4182_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6163_ (.A1(_3794_),
    .A2(_3796_),
    .A3(_1319_),
    .A4(_1179_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6164_ (.A1(_1182_),
    .A2(_1185_),
    .B(_1320_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6165_ (.A1(_0473_),
    .A2(\C[3][11] ),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _6166_ (.A1(_1184_),
    .A2(_4079_),
    .A3(_4176_),
    .A4(_1322_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _6167_ (.A1(_3961_),
    .A2(_4079_),
    .A3(_4093_),
    .B1(_1322_),
    .B2(_4088_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6168_ (.A1(_1323_),
    .A2(_1324_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6169_ (.A1(_3961_),
    .A2(_1020_),
    .A3(_4096_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6170_ (.A1(_1321_),
    .A2(_1325_),
    .A3(_1326_),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6171_ (.A1(_1318_),
    .A2(_1327_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6172_ (.A1(_1315_),
    .A2(_1328_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6173_ (.A1(_1311_),
    .A2(_1329_),
    .Z(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6174_ (.A1(_1307_),
    .A2(_1330_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6175_ (.A1(_1305_),
    .A2(_1331_),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6176_ (.A1(_1288_),
    .A2(_1291_),
    .A3(_1332_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6177_ (.A1(_1284_),
    .A2(_1333_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6178_ (.A1(_1282_),
    .A2(_1334_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6179_ (.A1(_1281_),
    .A2(_1335_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6180_ (.A1(_1194_),
    .A2(_1197_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6181_ (.A1(_1198_),
    .A2(_1203_),
    .B(_1337_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6182_ (.A1(_1336_),
    .A2(_1338_),
    .Z(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6183_ (.I(_1339_),
    .Z(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6184_ (.I(_1223_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6185_ (.A1(_1216_),
    .A2(_1340_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6186_ (.A1(_1061_),
    .A2(_1224_),
    .B(_1341_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6187_ (.A1(_1227_),
    .A2(_1268_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6188_ (.I(_1269_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6189_ (.A1(_1225_),
    .A2(_1344_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6190_ (.A1(_1343_),
    .A2(_1345_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6191_ (.A1(_1232_),
    .A2(_1236_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6192_ (.A1(_1228_),
    .A2(_1237_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6193_ (.A1(_1347_),
    .A2(_1348_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6194_ (.I(_0687_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6195_ (.A1(_0030_),
    .A2(_0054_),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6196_ (.A1(_0054_),
    .A2(_1234_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6197_ (.A1(_1234_),
    .A2(_1350_),
    .B(_1351_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6198_ (.I(_1352_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6199_ (.A1(_1221_),
    .A2(_1349_),
    .A3(_1353_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6200_ (.A1(_1242_),
    .A2(_1266_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6201_ (.A1(_1239_),
    .A2(_1267_),
    .B(_1355_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6202_ (.I(_1233_),
    .Z(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6203_ (.A1(_1262_),
    .A2(_1263_),
    .B(_1230_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6204_ (.A1(_1357_),
    .A2(_1358_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6205_ (.I(_1359_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6206_ (.A1(_1245_),
    .A2(_1258_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6207_ (.A1(_1259_),
    .A2(_1265_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6208_ (.A1(_1361_),
    .A2(_1362_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6209_ (.A1(_1253_),
    .A2(_1256_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6210_ (.A1(_1254_),
    .A2(_1255_),
    .B(_1364_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6211_ (.I(_1249_),
    .Z(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6212_ (.A1(_1366_),
    .A2(_1250_),
    .B(_1246_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6213_ (.A1(_1246_),
    .A2(_1366_),
    .A3(_1250_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6214_ (.A1(_1367_),
    .A2(_1257_),
    .B(_1368_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6215_ (.A1(_0981_),
    .A2(_0711_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6216_ (.I(_3972_),
    .Z(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6217_ (.I(_1371_),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6218_ (.A1(_1372_),
    .A2(\C[2][12] ),
    .A3(_0469_),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6219_ (.I(_1247_),
    .Z(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6220_ (.A1(_1374_),
    .A2(\C[2][12] ),
    .A3(\B[2][7] ),
    .A4(_0981_),
    .Z(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6221_ (.A1(_1370_),
    .A2(_1373_),
    .B(_1375_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6222_ (.A1(_1366_),
    .A2(_1376_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6223_ (.I(_1377_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6224_ (.A1(_1037_),
    .A2(_0037_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6225_ (.I(_0716_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6226_ (.A1(_4173_),
    .A2(_0039_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6227_ (.I(_0718_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6228_ (.A1(_4161_),
    .A2(_0038_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6229_ (.A1(_1379_),
    .A2(_1380_),
    .A3(_1381_),
    .Z(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6230_ (.A1(_1369_),
    .A2(_1378_),
    .A3(_1382_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6231_ (.A1(_1365_),
    .A2(_1383_),
    .Z(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6232_ (.A1(_1363_),
    .A2(_1384_),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6233_ (.A1(_1356_),
    .A2(_1360_),
    .A3(_1385_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6234_ (.A1(_1354_),
    .A2(_1386_),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6235_ (.A1(_1342_),
    .A2(_1346_),
    .A3(_1387_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6236_ (.A1(_1213_),
    .A2(_1270_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6237_ (.A1(_1213_),
    .A2(_1270_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6238_ (.A1(_1210_),
    .A2(_1389_),
    .B(_1390_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6239_ (.A1(_1388_),
    .A2(_1391_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6240_ (.A1(_1120_),
    .A2(_1272_),
    .A3(_1273_),
    .Z(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6241_ (.A1(_1121_),
    .A2(_1124_),
    .B(_1393_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6242_ (.A1(_1275_),
    .A2(_1272_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6243_ (.A1(_1273_),
    .A2(_1395_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6244_ (.A1(_1394_),
    .A2(_1396_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6245_ (.A1(_1392_),
    .A2(_1397_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6246_ (.I(_1398_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6247_ (.A1(_1194_),
    .A2(_1197_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6248_ (.A1(_1199_),
    .A2(_1202_),
    .B(_1336_),
    .C(_1399_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6249_ (.A1(_0985_),
    .A2(_1127_),
    .B(_1193_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6250_ (.A1(_1280_),
    .A2(_1401_),
    .A3(_1335_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6251_ (.A1(_1280_),
    .A2(_1401_),
    .B(_1335_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6252_ (.A1(_1194_),
    .A2(_1197_),
    .A3(_1402_),
    .B(_1403_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6253_ (.A1(_1400_),
    .A2(_1404_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6254_ (.A1(_1147_),
    .A2(_1287_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6255_ (.A1(_1291_),
    .A2(_1332_),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6256_ (.A1(_1291_),
    .A2(_1332_),
    .Z(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6257_ (.A1(_1288_),
    .A2(_1407_),
    .B(_1408_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6258_ (.A1(_1294_),
    .A2(_1304_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6259_ (.A1(_1167_),
    .A2(_1188_),
    .Z(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6260_ (.A1(_1306_),
    .A2(_1411_),
    .B(_1330_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6261_ (.A1(_1305_),
    .A2(_1331_),
    .B(_1412_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6262_ (.A1(_1298_),
    .A2(_1302_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6263_ (.A1(_0060_),
    .A2(_3900_),
    .A3(_1303_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6264_ (.A1(_1414_),
    .A2(_1415_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6265_ (.A1(_0061_),
    .A2(_3646_),
    .A3(_1301_),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6266_ (.A1(_1296_),
    .A2(_1300_),
    .B(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6267_ (.I(_1295_),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6268_ (.A1(_3326_),
    .A2(_1419_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6269_ (.I(_3874_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6270_ (.A1(_0062_),
    .A2(_3905_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6271_ (.A1(_3883_),
    .A2(_3899_),
    .ZN(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6272_ (.A1(_1420_),
    .A2(_1421_),
    .A3(_1422_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6273_ (.A1(_1418_),
    .A2(_1423_),
    .Z(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6274_ (.A1(_1416_),
    .A2(_1424_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6275_ (.I(_1311_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6276_ (.A1(_1315_),
    .A2(_1328_),
    .Z(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6277_ (.A1(_1426_),
    .A2(_1329_),
    .B(_1427_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6278_ (.A1(_1316_),
    .A2(_1317_),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6279_ (.A1(_1323_),
    .A2(_1324_),
    .A3(_1326_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6280_ (.A1(_1323_),
    .A2(_1324_),
    .B(_1326_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6281_ (.A1(_1321_),
    .A2(_1430_),
    .A3(_1431_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6282_ (.A1(_1318_),
    .A2(_1327_),
    .B(_1432_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6283_ (.A1(_0045_),
    .A2(_1037_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6284_ (.A1(_1184_),
    .A2(_4080_),
    .A3(_4176_),
    .A4(_1322_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6285_ (.A1(_1324_),
    .A2(_1326_),
    .B(_1435_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6286_ (.A1(_0456_),
    .A2(\C[3][12] ),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _6287_ (.A1(_4066_),
    .A2(_0755_),
    .A3(_4179_),
    .A4(_1437_),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6288_ (.A1(_3993_),
    .A2(_1020_),
    .A3(_4176_),
    .B1(_1437_),
    .B2(_4088_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6289_ (.A1(_1438_),
    .A2(_1439_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6290_ (.A1(_0335_),
    .A2(_3981_),
    .A3(_0337_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6291_ (.A1(_1436_),
    .A2(_1440_),
    .A3(_1441_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6292_ (.A1(_1434_),
    .A2(_1442_),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6293_ (.A1(_1433_),
    .A2(_1443_),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6294_ (.A1(_1429_),
    .A2(_1444_),
    .Z(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6295_ (.A1(_1428_),
    .A2(_1445_),
    .Z(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6296_ (.A1(_1425_),
    .A2(_1446_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6297_ (.A1(_1413_),
    .A2(_1447_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6298_ (.A1(_1410_),
    .A2(_1448_),
    .Z(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6299_ (.A1(_1409_),
    .A2(_1449_),
    .Z(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6300_ (.A1(_1406_),
    .A2(_1450_),
    .Z(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6301_ (.I(_1284_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6302_ (.A1(_1452_),
    .A2(_1333_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6303_ (.A1(_1282_),
    .A2(_1334_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6304_ (.A1(_1453_),
    .A2(_1454_),
    .Z(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6305_ (.A1(_1451_),
    .A2(_1455_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6306_ (.A1(_1405_),
    .A2(_1456_),
    .Z(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6307_ (.I(_1457_),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6308_ (.A1(_1346_),
    .A2(_1387_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6309_ (.A1(_1346_),
    .A2(_1387_),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6310_ (.A1(_1342_),
    .A2(_1458_),
    .A3(_1459_),
    .ZN(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6311_ (.A1(_1458_),
    .A2(_1460_),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6312_ (.A1(_1349_),
    .A2(_1353_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6313_ (.A1(_1349_),
    .A2(_1353_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6314_ (.A1(_1221_),
    .A2(_1462_),
    .B(_1463_),
    .ZN(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6315_ (.A1(_1359_),
    .A2(_1385_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6316_ (.A1(_1356_),
    .A2(_1465_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6317_ (.A1(_1354_),
    .A2(_1386_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6318_ (.A1(_1466_),
    .A2(_1467_),
    .ZN(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6319_ (.A1(_0031_),
    .A2(_0054_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6320_ (.A1(_1357_),
    .A2(_1358_),
    .B(_1469_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6321_ (.A1(_0327_),
    .A2(_1357_),
    .A3(_1358_),
    .B(_1470_),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6322_ (.A1(_1351_),
    .A2(_1471_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6323_ (.A1(_1380_),
    .A2(_1381_),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6324_ (.A1(_1380_),
    .A2(_1381_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6325_ (.A1(_1379_),
    .A2(_1473_),
    .B(_1474_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6326_ (.A1(_1378_),
    .A2(_1382_),
    .Z(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6327_ (.A1(_1366_),
    .A2(_1376_),
    .B(_1476_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6328_ (.A1(_3636_),
    .A2(_0711_),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6329_ (.I(_1374_),
    .Z(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6330_ (.A1(_1479_),
    .A2(\C[2][13] ),
    .A3(_0469_),
    .ZN(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6331_ (.A1(_1374_),
    .A2(\C[2][13] ),
    .A3(\B[2][7] ),
    .A4(_3625_),
    .Z(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6332_ (.A1(_1478_),
    .A2(_1480_),
    .B(_1481_),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6333_ (.A1(_1375_),
    .A2(_1482_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6334_ (.I(_1483_),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6335_ (.A1(_4161_),
    .A2(_0039_),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6336_ (.A1(_1038_),
    .A2(_0038_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6337_ (.A1(_1485_),
    .A2(_1486_),
    .Z(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6338_ (.A1(_1484_),
    .A2(_1487_),
    .Z(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6339_ (.A1(_1477_),
    .A2(_1488_),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6340_ (.A1(_1475_),
    .A2(_1489_),
    .Z(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6341_ (.A1(_1378_),
    .A2(_1382_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6342_ (.A1(_1369_),
    .A2(_1476_),
    .A3(_1491_),
    .B1(_1383_),
    .B2(_1365_),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6343_ (.A1(_1490_),
    .A2(_1492_),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6344_ (.A1(_1361_),
    .A2(_1362_),
    .B(_1384_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6345_ (.A1(_1360_),
    .A2(_1385_),
    .B(_1494_),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6346_ (.A1(_1493_),
    .A2(_1495_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6347_ (.A1(_1472_),
    .A2(_1496_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6348_ (.A1(_1468_),
    .A2(_1497_),
    .ZN(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6349_ (.A1(_1464_),
    .A2(_1498_),
    .Z(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6350_ (.A1(_1388_),
    .A2(_1391_),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6351_ (.A1(_1394_),
    .A2(_1396_),
    .B(_1392_),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6352_ (.A1(_1500_),
    .A2(_1501_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6353_ (.A1(_1461_),
    .A2(_1499_),
    .A3(_1502_),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6354_ (.I(_1503_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6355_ (.I(_1449_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6356_ (.A1(_1409_),
    .A2(_1504_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6357_ (.A1(_1406_),
    .A2(_1450_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6358_ (.A1(_1413_),
    .A2(_1447_),
    .Z(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6359_ (.A1(_1410_),
    .A2(_1448_),
    .B(_1507_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6360_ (.A1(_1416_),
    .A2(_1424_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6361_ (.A1(_1428_),
    .A2(_1445_),
    .Z(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6362_ (.A1(_1425_),
    .A2(_1446_),
    .B(_1510_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6363_ (.A1(_1418_),
    .A2(_1423_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6364_ (.I(_1421_),
    .Z(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6365_ (.A1(_3900_),
    .A2(_1419_),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6366_ (.A1(_1513_),
    .A2(_1514_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6367_ (.I(_1419_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6368_ (.A1(_0062_),
    .A2(_3900_),
    .B1(_3646_),
    .B2(_0063_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6369_ (.A1(_1515_),
    .A2(_1516_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6370_ (.A1(_3646_),
    .A2(_0063_),
    .ZN(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6371_ (.A1(_1420_),
    .A2(_1513_),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6372_ (.A1(_1300_),
    .A2(_1518_),
    .B1(_1422_),
    .B2(_1519_),
    .ZN(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6373_ (.A1(_1517_),
    .A2(_1520_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6374_ (.A1(_1512_),
    .A2(_1521_),
    .ZN(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6375_ (.A1(_1440_),
    .A2(_1441_),
    .Z(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6376_ (.A1(_1436_),
    .A2(_1523_),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6377_ (.A1(_3999_),
    .A2(_0023_),
    .A3(_1442_),
    .Z(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6378_ (.A1(_1524_),
    .A2(_1525_),
    .ZN(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6379_ (.A1(_3981_),
    .A2(_0339_),
    .A3(_1440_),
    .B(_1438_),
    .ZN(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6380_ (.I(_1372_),
    .Z(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6381_ (.I(_4085_),
    .Z(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6382_ (.I(_1529_),
    .Z(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6383_ (.A1(_4070_),
    .A2(_1530_),
    .ZN(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6384_ (.I(_1531_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6385_ (.A1(_1528_),
    .A2(\C[3][13] ),
    .A3(\A[2][6] ),
    .A4(_0047_),
    .ZN(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6386_ (.I(_1531_),
    .Z(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6387_ (.I(_0795_),
    .Z(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6388_ (.A1(_1479_),
    .A2(\C[3][13] ),
    .A3(_1534_),
    .ZN(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6389_ (.A1(_0337_),
    .A2(_1533_),
    .B(_1535_),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6390_ (.A1(_1532_),
    .A2(_1536_),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6391_ (.I(_3969_),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6392_ (.A1(_1538_),
    .A2(_0023_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6393_ (.A1(_1537_),
    .A2(_1539_),
    .Z(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6394_ (.A1(_1527_),
    .A2(_1540_),
    .Z(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6395_ (.I(_1541_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6396_ (.A1(_1526_),
    .A2(_1542_),
    .Z(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6397_ (.A1(_1433_),
    .A2(_1443_),
    .ZN(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6398_ (.A1(_1429_),
    .A2(_1444_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6399_ (.A1(_1544_),
    .A2(_1545_),
    .ZN(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6400_ (.A1(_1543_),
    .A2(_1546_),
    .Z(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6401_ (.A1(_1522_),
    .A2(_1547_),
    .Z(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6402_ (.A1(_1511_),
    .A2(_1548_),
    .Z(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6403_ (.A1(_1509_),
    .A2(_1549_),
    .Z(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6404_ (.A1(_1508_),
    .A2(_1550_),
    .Z(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6405_ (.A1(_1505_),
    .A2(_1506_),
    .B(_1551_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6406_ (.A1(_1505_),
    .A2(_1506_),
    .A3(_1551_),
    .Z(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6407_ (.A1(_1552_),
    .A2(_1553_),
    .Z(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6408_ (.A1(_1453_),
    .A2(_1454_),
    .B(_1451_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6409_ (.A1(_1405_),
    .A2(_1456_),
    .B(_1555_),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6410_ (.A1(_1554_),
    .A2(_1556_),
    .Z(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6411_ (.I(_1557_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6412_ (.A1(_1468_),
    .A2(_1497_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6413_ (.I(_1464_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6414_ (.A1(_1559_),
    .A2(_1498_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6415_ (.A1(_0327_),
    .A2(_1357_),
    .A3(_1358_),
    .B1(_1471_),
    .B2(_1351_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6416_ (.A1(_1493_),
    .A2(_1495_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6417_ (.A1(_1472_),
    .A2(_1496_),
    .B(_1562_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6418_ (.A1(_1490_),
    .A2(_1492_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6419_ (.I(_1488_),
    .ZN(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6420_ (.A1(_1477_),
    .A2(_1565_),
    .ZN(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6421_ (.A1(_1475_),
    .A2(_1489_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6422_ (.A1(_1566_),
    .A2(_1567_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6423_ (.A1(_1485_),
    .A2(_1486_),
    .Z(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6424_ (.A1(_1528_),
    .A2(\C[2][14] ),
    .A3(\B[2][7] ),
    .A4(_3898_),
    .Z(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6425_ (.A1(\C[2][14] ),
    .A2(_0185_),
    .B1(_1094_),
    .B2(_3898_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6426_ (.A1(_1570_),
    .A2(_1571_),
    .ZN(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6427_ (.A1(_1481_),
    .A2(_1572_),
    .ZN(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6428_ (.A1(_1038_),
    .A2(_0039_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6429_ (.A1(_1573_),
    .A2(_1574_),
    .ZN(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6430_ (.A1(_1375_),
    .A2(_1482_),
    .B1(_1484_),
    .B2(_1487_),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6431_ (.A1(_1575_),
    .A2(_1576_),
    .ZN(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6432_ (.A1(_1569_),
    .A2(_1577_),
    .ZN(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6433_ (.A1(_1568_),
    .A2(_1578_),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6434_ (.A1(_1564_),
    .A2(_1579_),
    .Z(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6435_ (.A1(_1563_),
    .A2(_1580_),
    .Z(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6436_ (.A1(_1561_),
    .A2(_1581_),
    .Z(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6437_ (.A1(_1558_),
    .A2(_1560_),
    .B(_1582_),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6438_ (.A1(_1558_),
    .A2(_1560_),
    .A3(_1582_),
    .Z(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6439_ (.A1(_1583_),
    .A2(_1584_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6440_ (.A1(_1458_),
    .A2(_1460_),
    .B(_1499_),
    .ZN(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6441_ (.A1(_1458_),
    .A2(_1460_),
    .A3(_1499_),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6442_ (.A1(_1500_),
    .A2(_1501_),
    .A3(_1586_),
    .B(_1587_),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6443_ (.A1(_1585_),
    .A2(_1588_),
    .Z(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6444_ (.I(_1589_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6445_ (.A1(_1508_),
    .A2(_1550_),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6446_ (.A1(_1512_),
    .A2(_1521_),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6447_ (.A1(_1517_),
    .A2(_1520_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6448_ (.A1(_0031_),
    .A2(_0063_),
    .A3(_1513_),
    .ZN(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6449_ (.A1(_1592_),
    .A2(_1593_),
    .ZN(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6450_ (.A1(_1537_),
    .A2(_1539_),
    .B(_1532_),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6451_ (.A1(_4152_),
    .A2(_1533_),
    .ZN(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6452_ (.I(_1528_),
    .Z(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6453_ (.I(_1597_),
    .Z(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6454_ (.A1(_1598_),
    .A2(\C[3][14] ),
    .A3(_1534_),
    .Z(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6455_ (.A1(_1598_),
    .A2(\C[3][14] ),
    .A3(_1596_),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6456_ (.A1(_1596_),
    .A2(_1599_),
    .B(_1600_),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6457_ (.I(_1601_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6458_ (.A1(_1595_),
    .A2(_1602_),
    .Z(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6459_ (.A1(_1527_),
    .A2(_1540_),
    .Z(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6460_ (.A1(_1526_),
    .A2(_1542_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6461_ (.A1(_1604_),
    .A2(_1605_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6462_ (.A1(_1603_),
    .A2(_1606_),
    .Z(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6463_ (.A1(_1594_),
    .A2(_1607_),
    .Z(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6464_ (.A1(_1544_),
    .A2(_1545_),
    .B(_1543_),
    .ZN(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6465_ (.A1(_1522_),
    .A2(_1547_),
    .B(_1609_),
    .ZN(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6466_ (.A1(_1608_),
    .A2(_1610_),
    .ZN(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6467_ (.A1(_1591_),
    .A2(_1611_),
    .Z(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6468_ (.I(_1511_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6469_ (.A1(_1613_),
    .A2(_1548_),
    .ZN(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6470_ (.A1(_1509_),
    .A2(_1549_),
    .B(_1614_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6471_ (.A1(_1612_),
    .A2(_1615_),
    .Z(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6472_ (.A1(_1590_),
    .A2(_1616_),
    .ZN(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6473_ (.A1(_1555_),
    .A2(_1552_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6474_ (.A1(_1553_),
    .A2(_1618_),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6475_ (.A1(_1451_),
    .A2(_1455_),
    .Z(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6476_ (.A1(_1400_),
    .A2(_1404_),
    .B(_1620_),
    .C(_1554_),
    .ZN(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6477_ (.A1(_1619_),
    .A2(_1621_),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6478_ (.A1(_1617_),
    .A2(_1622_),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6479_ (.I(_1623_),
    .Z(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6480_ (.A1(_1563_),
    .A2(_1580_),
    .ZN(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6481_ (.A1(_1561_),
    .A2(_1581_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6482_ (.A1(_1568_),
    .A2(_1578_),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6483_ (.A1(_1564_),
    .A2(_1579_),
    .ZN(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6484_ (.I(_0947_),
    .Z(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6485_ (.A1(\C[2][15] ),
    .A2(_1628_),
    .Z(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6486_ (.I(_1534_),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6487_ (.A1(\C[2][15] ),
    .A2(_1630_),
    .A3(_1570_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6488_ (.A1(_1570_),
    .A2(_1629_),
    .B(_1631_),
    .ZN(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6489_ (.A1(_1573_),
    .A2(_1574_),
    .ZN(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6490_ (.A1(_1481_),
    .A2(_1572_),
    .B(_1633_),
    .ZN(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6491_ (.A1(_1575_),
    .A2(_1576_),
    .ZN(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6492_ (.A1(_1569_),
    .A2(_1577_),
    .ZN(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6493_ (.A1(_1635_),
    .A2(_1636_),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6494_ (.A1(_1632_),
    .A2(_1634_),
    .A3(_1637_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6495_ (.A1(_1626_),
    .A2(_1627_),
    .B(_1638_),
    .ZN(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6496_ (.A1(_1626_),
    .A2(_1627_),
    .A3(_1638_),
    .Z(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6497_ (.A1(_1639_),
    .A2(_1640_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6498_ (.A1(_1624_),
    .A2(_1625_),
    .B(_1641_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6499_ (.A1(_1624_),
    .A2(_1625_),
    .A3(_1641_),
    .Z(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6500_ (.A1(_1642_),
    .A2(_1643_),
    .ZN(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6501_ (.A1(_1585_),
    .A2(_1588_),
    .B(_1583_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6502_ (.A1(_1644_),
    .A2(_1645_),
    .Z(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6503_ (.I(_1646_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6504_ (.A1(_1590_),
    .A2(_1616_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6505_ (.A1(_1619_),
    .A2(_1621_),
    .B(_1617_),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6506_ (.I(_1612_),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6507_ (.A1(_1649_),
    .A2(_1615_),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6508_ (.A1(_1592_),
    .A2(_1593_),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6509_ (.A1(_1608_),
    .A2(_1610_),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6510_ (.A1(_1512_),
    .A2(_1521_),
    .A3(_1611_),
    .B(_1652_),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6511_ (.A1(_1605_),
    .A2(_1603_),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6512_ (.A1(_1594_),
    .A2(_1607_),
    .B(_1654_),
    .ZN(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6513_ (.A1(_1604_),
    .A2(_1603_),
    .Z(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6514_ (.A1(_1595_),
    .A2(_1602_),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6515_ (.A1(_1600_),
    .A2(_1657_),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6516_ (.A1(\C[3][15] ),
    .A2(_0947_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6517_ (.A1(_1658_),
    .A2(_1659_),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6518_ (.A1(_1656_),
    .A2(_1660_),
    .ZN(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6519_ (.A1(_1515_),
    .A2(_1661_),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6520_ (.A1(_1655_),
    .A2(_1662_),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6521_ (.A1(_1651_),
    .A2(_1653_),
    .A3(_1663_),
    .Z(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6522_ (.A1(_1650_),
    .A2(_1664_),
    .Z(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6523_ (.A1(_1647_),
    .A2(_1648_),
    .A3(_1665_),
    .Z(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6524_ (.A1(_1647_),
    .A2(_1648_),
    .B(_1665_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6525_ (.A1(_1666_),
    .A2(_1667_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6526_ (.A1(_1585_),
    .A2(_1642_),
    .A3(_1643_),
    .Z(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6527_ (.I(_1642_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6528_ (.A1(_1583_),
    .A2(_1643_),
    .B1(_1668_),
    .B2(_1588_),
    .C(_1669_),
    .ZN(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6529_ (.I(\C[2][16] ),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6530_ (.I(_4087_),
    .Z(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6531_ (.I(_1672_),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6532_ (.A1(_3434_),
    .A2(_1671_),
    .A3(_1673_),
    .B(_1631_),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6533_ (.A1(_3434_),
    .A2(_1671_),
    .A3(_1631_),
    .B(_1674_),
    .ZN(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6534_ (.A1(_1632_),
    .A2(_1634_),
    .Z(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6535_ (.A1(_1632_),
    .A2(_1634_),
    .Z(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6536_ (.A1(_1676_),
    .A2(_1637_),
    .B(_1677_),
    .ZN(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6537_ (.A1(_1639_),
    .A2(_1675_),
    .A3(_1678_),
    .Z(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6538_ (.A1(_1670_),
    .A2(_1679_),
    .Z(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6539_ (.I(_1680_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6540_ (.A1(_1619_),
    .A2(_1621_),
    .B(_1665_),
    .C(_1617_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6541_ (.A1(_1590_),
    .A2(_1616_),
    .B(_1650_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6542_ (.A1(_1664_),
    .A2(_1682_),
    .Z(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6543_ (.A1(_1513_),
    .A2(_1514_),
    .A3(_1661_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6544_ (.A1(_1657_),
    .A2(_1659_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6545_ (.A1(_1656_),
    .A2(_1660_),
    .B(_1684_),
    .C(_1685_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6546_ (.A1(\C[3][15] ),
    .A2(_1596_),
    .A3(_1599_),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6547_ (.I(_1598_),
    .Z(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6548_ (.A1(_1688_),
    .A2(\C[3][16] ),
    .Z(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6549_ (.A1(\C[3][16] ),
    .A2(_1628_),
    .A3(_1687_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6550_ (.A1(_1687_),
    .A2(_1689_),
    .B(_1690_),
    .ZN(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6551_ (.A1(_1651_),
    .A2(_1663_),
    .Z(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6552_ (.A1(_1651_),
    .A2(_1663_),
    .Z(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6553_ (.A1(_1655_),
    .A2(_1662_),
    .B1(_1692_),
    .B2(_1653_),
    .C(_1693_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6554_ (.A1(_1686_),
    .A2(_1691_),
    .A3(_1694_),
    .ZN(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6555_ (.A1(_1681_),
    .A2(_1683_),
    .A3(_1695_),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6556_ (.A1(_1681_),
    .A2(_1683_),
    .B(_1695_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6557_ (.A1(_1696_),
    .A2(_1697_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _6558_ (.A1(_3779_),
    .A2(_3445_),
    .A3(_3782_),
    .ZN(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6559_ (.A1(_2481_),
    .A2(_3746_),
    .A3(_3747_),
    .A4(_2287_),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _6560_ (.A1(_3380_),
    .A2(_1698_),
    .B1(_1699_),
    .B2(\A[1][0] ),
    .C(_3759_),
    .ZN(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6561_ (.I(_1700_),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6562_ (.I(_1701_),
    .Z(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6563_ (.I(_1702_),
    .Z(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6564_ (.I(_1703_),
    .Z(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6565_ (.A1(_0208_),
    .A2(_1704_),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6566_ (.I(_3809_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6567_ (.A1(_2244_),
    .A2(_2265_),
    .A3(_2383_),
    .ZN(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6568_ (.I(_1706_),
    .Z(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6569_ (.A1(_3358_),
    .A2(_3369_),
    .A3(_1707_),
    .ZN(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _6570_ (.A1(net3),
    .A2(net2),
    .A3(net4),
    .Z(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6571_ (.I(_1709_),
    .Z(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6572_ (.I(\A[0][0] ),
    .ZN(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6573_ (.A1(_3531_),
    .A2(_1710_),
    .B(_1711_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _6574_ (.A1(_1708_),
    .A2(_1712_),
    .Z(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6575_ (.I(_1713_),
    .Z(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6576_ (.I(_1714_),
    .Z(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6577_ (.I(_1715_),
    .Z(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6578_ (.A1(_0040_),
    .A2(_1716_),
    .ZN(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6579_ (.A1(_1688_),
    .A2(\C[1][0] ),
    .A3(_1630_),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6580_ (.A1(_1479_),
    .A2(\C[1][0] ),
    .A3(_0040_),
    .A4(_1715_),
    .Z(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6581_ (.A1(_1717_),
    .A2(_1718_),
    .B(_1719_),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6582_ (.A1(_1705_),
    .A2(_1720_),
    .Z(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6583_ (.I(_1721_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6584_ (.A1(_1705_),
    .A2(_1720_),
    .Z(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6585_ (.I(\B[1][1] ),
    .Z(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6586_ (.A1(_3759_),
    .A2(_1708_),
    .A3(_1712_),
    .ZN(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6587_ (.I(_1724_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6588_ (.I(_1725_),
    .Z(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _6589_ (.A1(_1371_),
    .A2(\C[1][1] ),
    .A3(_1723_),
    .A4(_1726_),
    .Z(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6590_ (.I(_1726_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6591_ (.A1(_1371_),
    .A2(\C[1][1] ),
    .A3(_0468_),
    .Z(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6592_ (.A1(_4157_),
    .A2(_0000_),
    .B(_1728_),
    .ZN(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6593_ (.A1(_1727_),
    .A2(_1729_),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6594_ (.I(_1709_),
    .Z(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _6595_ (.A1(_3037_),
    .A2(_1731_),
    .B(\A[0][1] ),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6596_ (.I(_1707_),
    .Z(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6597_ (.A1(_3078_),
    .A2(_1733_),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6598_ (.A1(_1732_),
    .A2(_1734_),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6599_ (.I(_1735_),
    .Z(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6600_ (.A1(_0040_),
    .A2(_1736_),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6601_ (.A1(_1719_),
    .A2(_1730_),
    .A3(_1737_),
    .Z(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6602_ (.I(_1700_),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6603_ (.I(_1739_),
    .Z(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6604_ (.A1(_0211_),
    .A2(_1740_),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _6605_ (.A1(_3746_),
    .A2(_3748_),
    .A3(_2394_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _6606_ (.A1(_3358_),
    .A2(_3779_),
    .A3(_2373_),
    .A4(_2567_),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6607_ (.A1(_3797_),
    .A2(_1742_),
    .B1(_1743_),
    .B2(\A[1][1] ),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6608_ (.A1(_3792_),
    .A2(_1744_),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6609_ (.I(_1745_),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6610_ (.I(_1746_),
    .Z(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6611_ (.I(_1747_),
    .Z(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6612_ (.A1(_3488_),
    .A2(_1748_),
    .ZN(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6613_ (.A1(_1741_),
    .A2(_1749_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6614_ (.A1(_1738_),
    .A2(_1750_),
    .Z(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6615_ (.A1(_1722_),
    .A2(_1751_),
    .Z(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6616_ (.I(_1752_),
    .Z(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6617_ (.I(_2867_),
    .Z(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6618_ (.A1(_2816_),
    .A2(_1742_),
    .B1(_1743_),
    .B2(\A[1][2] ),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6619_ (.I(_1754_),
    .Z(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6620_ (.A1(_1753_),
    .A2(_1755_),
    .Z(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6621_ (.I(_1756_),
    .Z(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6622_ (.I(_1757_),
    .Z(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6623_ (.I(_1758_),
    .Z(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6624_ (.A1(_3904_),
    .A2(_1740_),
    .A3(_1749_),
    .A4(_1759_),
    .Z(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6625_ (.I(_1745_),
    .ZN(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6626_ (.I(_1761_),
    .Z(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6627_ (.I(_1762_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6628_ (.A1(_0208_),
    .A2(_1759_),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6629_ (.A1(_0211_),
    .A2(_0009_),
    .B(_1763_),
    .ZN(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6630_ (.I(_1756_),
    .ZN(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6631_ (.A1(_4116_),
    .A2(_1703_),
    .A3(_1749_),
    .A4(_1765_),
    .Z(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6632_ (.A1(_1760_),
    .A2(_1764_),
    .A3(_1766_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6633_ (.I(_2427_),
    .Z(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6634_ (.A1(_1768_),
    .A2(_1702_),
    .ZN(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6635_ (.I(_1724_),
    .Z(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6636_ (.I(_1770_),
    .Z(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6637_ (.I(_1771_),
    .Z(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6638_ (.A1(_3786_),
    .A2(_1772_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6639_ (.A1(_1769_),
    .A2(_1773_),
    .Z(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6640_ (.I(\A[0][1] ),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6641_ (.A1(_3185_),
    .A2(_1733_),
    .B(_1775_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6642_ (.I(_1710_),
    .Z(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6643_ (.A1(_3196_),
    .A2(_1777_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6644_ (.A1(_1776_),
    .A2(_1778_),
    .B(_3760_),
    .ZN(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6645_ (.I(_1779_),
    .ZN(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6646_ (.I(_1780_),
    .Z(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6647_ (.A1(_0457_),
    .A2(\C[1][2] ),
    .A3(_1723_),
    .A4(_1781_),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6648_ (.I(net38),
    .Z(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6649_ (.A1(_3972_),
    .A2(\C[1][2] ),
    .A3(_3975_),
    .Z(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6650_ (.A1(_4157_),
    .A2(_1783_),
    .B(_1784_),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6651_ (.A1(_1782_),
    .A2(_1785_),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6652_ (.I(\A[0][2] ),
    .ZN(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6653_ (.A1(_3402_),
    .A2(_1707_),
    .B(_1787_),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6654_ (.A1(_2341_),
    .A2(_1710_),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6655_ (.A1(_1788_),
    .A2(_1789_),
    .B(_3759_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6656_ (.I(net34),
    .Z(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6657_ (.A1(_0179_),
    .A2(_1791_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6658_ (.A1(_1727_),
    .A2(_1786_),
    .A3(_1792_),
    .Z(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6659_ (.A1(_1727_),
    .A2(_1729_),
    .B(_1737_),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6660_ (.A1(_1727_),
    .A2(_1729_),
    .A3(_1737_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6661_ (.A1(_1719_),
    .A2(_1794_),
    .B(_1795_),
    .ZN(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6662_ (.A1(_1793_),
    .A2(_1796_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6663_ (.A1(_1774_),
    .A2(_1797_),
    .Z(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6664_ (.A1(_1767_),
    .A2(_1798_),
    .Z(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6665_ (.I(_1799_),
    .ZN(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6666_ (.A1(_1738_),
    .A2(_1750_),
    .ZN(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6667_ (.A1(_1722_),
    .A2(_1751_),
    .B(_1801_),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6668_ (.A1(_1800_),
    .A2(_1802_),
    .Z(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6669_ (.I(_1803_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6670_ (.A1(_1722_),
    .A2(_1751_),
    .A3(_1799_),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6671_ (.A1(_1801_),
    .A2(_1799_),
    .ZN(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6672_ (.A1(_1767_),
    .A2(_1798_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6673_ (.I(_1765_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _6674_ (.A1(_2897_),
    .A2(_1742_),
    .B1(_1743_),
    .B2(\A[1][3] ),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6675_ (.A1(_3776_),
    .A2(_1807_),
    .Z(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6676_ (.I(_1808_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6677_ (.I(_1809_),
    .Z(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6678_ (.I(_1810_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6679_ (.I(_1811_),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6680_ (.A1(_0202_),
    .A2(_0010_),
    .B1(_1812_),
    .B2(_3510_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6681_ (.I(_1808_),
    .Z(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6682_ (.A1(_4116_),
    .A2(_0009_),
    .A3(_1763_),
    .A4(_1814_),
    .ZN(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6683_ (.A1(_0211_),
    .A2(_1748_),
    .A3(_1763_),
    .A4(_1812_),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6684_ (.A1(_1815_),
    .A2(_1816_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6685_ (.A1(_1813_),
    .A2(_1817_),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6686_ (.I(_1795_),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6687_ (.A1(_1719_),
    .A2(_1819_),
    .A3(_1794_),
    .A4(_1793_),
    .Z(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6688_ (.A1(_1774_),
    .A2(_1797_),
    .B(_1820_),
    .ZN(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6689_ (.A1(_1769_),
    .A2(_1773_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6690_ (.I(_1700_),
    .Z(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6691_ (.A1(_4200_),
    .A2(_1823_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6692_ (.A1(_1768_),
    .A2(_1747_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6693_ (.I(_1780_),
    .Z(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6694_ (.I(_1826_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6695_ (.A1(_4215_),
    .A2(_0001_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6696_ (.A1(_1824_),
    .A2(_1825_),
    .A3(_1827_),
    .Z(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6697_ (.A1(_1822_),
    .A2(_1828_),
    .Z(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6698_ (.I(_1829_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6699_ (.A1(_1795_),
    .A2(_1793_),
    .ZN(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6700_ (.A1(_3962_),
    .A2(_1772_),
    .ZN(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6701_ (.A1(_1374_),
    .A2(\C[1][1] ),
    .A3(_1723_),
    .A4(_0000_),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6702_ (.A1(_1782_),
    .A2(_1785_),
    .B(_1833_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6703_ (.A1(_1833_),
    .A2(_1782_),
    .A3(_1785_),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6704_ (.A1(_1834_),
    .A2(_1792_),
    .B(_1835_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6705_ (.A1(_1247_),
    .A2(\C[1][2] ),
    .A3(_1723_),
    .A4(_1781_),
    .ZN(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6706_ (.I(_3766_),
    .Z(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6707_ (.I(_1790_),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6708_ (.I(_1839_),
    .Z(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6709_ (.I(_1840_),
    .Z(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6710_ (.A1(_0513_),
    .A2(\C[1][3] ),
    .Z(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6711_ (.A1(_1838_),
    .A2(_1841_),
    .A3(_1842_),
    .Z(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6712_ (.A1(_4009_),
    .A2(_1841_),
    .B1(_1842_),
    .B2(_3975_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6713_ (.A1(_1843_),
    .A2(_1844_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6714_ (.A1(_2492_),
    .A2(_1731_),
    .B(\A[0][3] ),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6715_ (.I(_1846_),
    .Z(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6716_ (.I(_1706_),
    .Z(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6717_ (.A1(_2599_),
    .A2(_1848_),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6718_ (.I(_1849_),
    .Z(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6719_ (.A1(_1847_),
    .A2(_1850_),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6720_ (.A1(_4012_),
    .A2(_1851_),
    .Z(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6721_ (.A1(_1837_),
    .A2(_1845_),
    .A3(_1852_),
    .Z(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6722_ (.A1(_1836_),
    .A2(_1853_),
    .Z(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6723_ (.A1(_1831_),
    .A2(_1832_),
    .A3(_1854_),
    .Z(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _6724_ (.A1(_1821_),
    .A2(_1830_),
    .A3(_1855_),
    .Z(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6725_ (.A1(_1806_),
    .A2(_1818_),
    .A3(_1856_),
    .Z(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6726_ (.A1(_1760_),
    .A2(_1805_),
    .A3(_1857_),
    .Z(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6727_ (.A1(_1804_),
    .A2(_1858_),
    .Z(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6728_ (.I(_1859_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6729_ (.I(\A[1][4] ),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6730_ (.I(_1699_),
    .Z(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _6731_ (.A1(_1860_),
    .A2(_2674_),
    .A3(_1861_),
    .B1(_1698_),
    .B2(_3802_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6732_ (.I(_1862_),
    .Z(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6733_ (.I(_1863_),
    .Z(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6734_ (.I(_1864_),
    .Z(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6735_ (.I(_1865_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6736_ (.I(_1740_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6737_ (.A1(_0057_),
    .A2(_0008_),
    .A3(_1749_),
    .A4(_1759_),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6738_ (.A1(_1818_),
    .A2(_1856_),
    .Z(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6739_ (.A1(_1866_),
    .A2(_1867_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6740_ (.A1(_1760_),
    .A2(_1857_),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6741_ (.A1(_1722_),
    .A2(_1751_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _6742_ (.A1(_1805_),
    .A2(_1868_),
    .A3(_1869_),
    .B1(_1858_),
    .B2(_1870_),
    .B3(_1800_),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6743_ (.A1(_1866_),
    .A2(_1806_),
    .B(_1867_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6744_ (.A1(_1829_),
    .A2(_1855_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _6745_ (.A1(_1813_),
    .A2(_1817_),
    .A3(_1856_),
    .B1(_1873_),
    .B2(net36),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6746_ (.A1(_1832_),
    .A2(_1854_),
    .Z(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6747_ (.A1(_1832_),
    .A2(_1854_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6748_ (.A1(_1831_),
    .A2(_1875_),
    .A3(_1876_),
    .B1(_1855_),
    .B2(_1830_),
    .ZN(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6749_ (.A1(_4200_),
    .A2(_1746_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6750_ (.A1(_1824_),
    .A2(_1825_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6751_ (.A1(_1769_),
    .A2(_1878_),
    .B(_1879_),
    .C(_1827_),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6752_ (.A1(_2449_),
    .A2(_1765_),
    .ZN(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6753_ (.I(_1739_),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6754_ (.A1(_4202_),
    .A2(_1882_),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6755_ (.A1(_1878_),
    .A2(_1881_),
    .A3(_1883_),
    .Z(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6756_ (.A1(_3786_),
    .A2(_1791_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6757_ (.A1(_1884_),
    .A2(_1885_),
    .Z(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6758_ (.A1(_1880_),
    .A2(_1886_),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6759_ (.A1(_1836_),
    .A2(_1853_),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _6760_ (.A1(_3962_),
    .A2(_1772_),
    .A3(_1888_),
    .B1(_1853_),
    .B2(_1836_),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6761_ (.A1(_4076_),
    .A2(_0001_),
    .ZN(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6762_ (.A1(_1843_),
    .A2(_1844_),
    .B(_1837_),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6763_ (.A1(_1837_),
    .A2(_1843_),
    .A3(_1844_),
    .ZN(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6764_ (.A1(_1891_),
    .A2(_1852_),
    .B(_1892_),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6765_ (.I(_1840_),
    .Z(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6766_ (.A1(_3767_),
    .A2(_1894_),
    .A3(_1842_),
    .ZN(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6767_ (.A1(_3931_),
    .A2(_1725_),
    .ZN(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6768_ (.A1(_3542_),
    .A2(_1777_),
    .B(\A[0][4] ),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6769_ (.A1(_3819_),
    .A2(_1733_),
    .ZN(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6770_ (.A1(_1897_),
    .A2(_1898_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6771_ (.A1(_3832_),
    .A2(_1899_),
    .ZN(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6772_ (.A1(_1896_),
    .A2(_1900_),
    .Z(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6773_ (.A1(_1846_),
    .A2(_1849_),
    .B(_2674_),
    .ZN(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6774_ (.I(_1902_),
    .Z(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6775_ (.A1(_3971_),
    .A2(\C[1][4] ),
    .Z(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6776_ (.A1(_1838_),
    .A2(_1903_),
    .A3(_1904_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6777_ (.I(_1905_),
    .Z(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6778_ (.I(_1903_),
    .Z(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _6779_ (.A1(_3767_),
    .A2(_1907_),
    .B1(_1904_),
    .B2(_0476_),
    .ZN(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6780_ (.A1(_1906_),
    .A2(_1908_),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6781_ (.A1(_1895_),
    .A2(_1901_),
    .A3(_1909_),
    .Z(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6782_ (.A1(_1893_),
    .A2(_1910_),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6783_ (.A1(_1890_),
    .A2(_1911_),
    .Z(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6784_ (.A1(_1887_),
    .A2(_1889_),
    .A3(_1912_),
    .ZN(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6785_ (.I(_1812_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6786_ (.A1(_0202_),
    .A2(_1763_),
    .A3(_0011_),
    .ZN(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6787_ (.A1(_1822_),
    .A2(_1828_),
    .ZN(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6788_ (.A1(_3229_),
    .A2(_1811_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6789_ (.A1(_4113_),
    .A2(_1762_),
    .A3(_1824_),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6790_ (.A1(_1916_),
    .A2(_1917_),
    .Z(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6791_ (.A1(_3888_),
    .A2(_1865_),
    .ZN(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6792_ (.A1(_1918_),
    .A2(_1919_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6793_ (.A1(_1915_),
    .A2(_1920_),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6794_ (.A1(_1914_),
    .A2(_1921_),
    .Z(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6795_ (.A1(_1877_),
    .A2(_1913_),
    .A3(_1922_),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6796_ (.A1(_1815_),
    .A2(_1874_),
    .A3(_1923_),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6797_ (.A1(_1871_),
    .A2(_1872_),
    .A3(_1924_),
    .Z(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6798_ (.I(_1925_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6799_ (.I(\A[1][5] ),
    .ZN(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _6800_ (.A1(_1926_),
    .A2(_3775_),
    .A3(_1861_),
    .B1(_1698_),
    .B2(_3829_),
    .ZN(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6801_ (.I(_1927_),
    .Z(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6802_ (.I(_1928_),
    .Z(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6803_ (.I(_1929_),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6804_ (.I(_1930_),
    .Z(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6805_ (.I(_1931_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6806_ (.A1(_1872_),
    .A2(_1924_),
    .Z(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6807_ (.A1(_1872_),
    .A2(_1924_),
    .Z(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6808_ (.A1(_1871_),
    .A2(_1932_),
    .B(_1933_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6809_ (.A1(_1874_),
    .A2(_1923_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6810_ (.A1(net35),
    .A2(_1923_),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6811_ (.A1(_1815_),
    .A2(_1935_),
    .B(_1936_),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6812_ (.A1(_1915_),
    .A2(_1920_),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6813_ (.A1(_1914_),
    .A2(_1921_),
    .B(_1938_),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6814_ (.A1(_1877_),
    .A2(_1913_),
    .Z(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6815_ (.A1(_1877_),
    .A2(_1913_),
    .Z(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6816_ (.A1(_1940_),
    .A2(_1922_),
    .B(_1941_),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6817_ (.A1(_3889_),
    .A2(_0012_),
    .A3(_1918_),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6818_ (.A1(_1916_),
    .A2(_1917_),
    .B(_1943_),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6819_ (.A1(_1880_),
    .A2(_1886_),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6820_ (.A1(_4202_),
    .A2(_1740_),
    .B1(_1761_),
    .B2(_4195_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6821_ (.A1(_0980_),
    .A2(_1761_),
    .A3(_1824_),
    .ZN(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6822_ (.A1(_1881_),
    .A2(_1946_),
    .B(_1947_),
    .ZN(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6823_ (.I(_1864_),
    .Z(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6824_ (.A1(_3218_),
    .A2(_1949_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6825_ (.A1(_1948_),
    .A2(_1950_),
    .ZN(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6826_ (.I(_1930_),
    .Z(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6827_ (.A1(_3499_),
    .A2(_1952_),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6828_ (.A1(_1951_),
    .A2(_1953_),
    .Z(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6829_ (.A1(_1945_),
    .A2(_1954_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6830_ (.A1(_1944_),
    .A2(_1955_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6831_ (.A1(net39),
    .A2(_1912_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6832_ (.A1(net39),
    .A2(_1912_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6833_ (.A1(_1887_),
    .A2(_1957_),
    .B(_1958_),
    .ZN(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6834_ (.A1(_1884_),
    .A2(_1885_),
    .ZN(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6835_ (.A1(_3864_),
    .A2(_1882_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6836_ (.I(_1902_),
    .Z(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6837_ (.A1(_4007_),
    .A2(_1962_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6838_ (.A1(_1961_),
    .A2(_1963_),
    .Z(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6839_ (.A1(_3004_),
    .A2(_1747_),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6840_ (.A1(_2460_),
    .A2(_1811_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6841_ (.A1(_4200_),
    .A2(_1758_),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6842_ (.A1(_1965_),
    .A2(_1966_),
    .A3(_1967_),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6843_ (.A1(_1964_),
    .A2(_1968_),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6844_ (.A1(_1960_),
    .A2(_1969_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6845_ (.I(_1779_),
    .Z(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6846_ (.I(_1971_),
    .Z(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6847_ (.A1(_3962_),
    .A2(_1972_),
    .A3(_1911_),
    .B1(_1910_),
    .B2(_1893_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6848_ (.A1(_1896_),
    .A2(_1900_),
    .Z(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6849_ (.I(_1839_),
    .Z(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6850_ (.I(_1975_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6851_ (.A1(_4076_),
    .A2(_0002_),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6852_ (.A1(_1906_),
    .A2(_1908_),
    .B(_1895_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6853_ (.A1(_1895_),
    .A2(_1906_),
    .A3(_1908_),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6854_ (.A1(_1901_),
    .A2(_1977_),
    .B(_1978_),
    .ZN(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _6855_ (.I(_1971_),
    .Z(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6856_ (.A1(_2492_),
    .A2(_1731_),
    .B(\A[0][5] ),
    .ZN(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6857_ (.A1(_3260_),
    .A2(_1848_),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6858_ (.A1(_1981_),
    .A2(_1982_),
    .Z(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6859_ (.A1(_4001_),
    .A2(_4150_),
    .A3(_1980_),
    .A4(_1983_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6860_ (.I(_3931_),
    .Z(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6861_ (.A1(_1981_),
    .A2(_1982_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6862_ (.I(_1986_),
    .Z(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6863_ (.A1(_1985_),
    .A2(_1783_),
    .B1(_1987_),
    .B2(_4012_),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6864_ (.A1(_1984_),
    .A2(_1988_),
    .ZN(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6865_ (.A1(_3982_),
    .A2(\C[1][5] ),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6866_ (.A1(_3949_),
    .A2(_1724_),
    .A3(_1990_),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6867_ (.A1(_4087_),
    .A2(_1990_),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6868_ (.A1(_3957_),
    .A2(_1725_),
    .B(_1992_),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6869_ (.A1(_1991_),
    .A2(_1993_),
    .ZN(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6870_ (.I(\A[0][4] ),
    .ZN(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6871_ (.A1(_2330_),
    .A2(_1707_),
    .B(_1995_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6872_ (.A1(_3802_),
    .A2(_1710_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6873_ (.A1(_1996_),
    .A2(_1997_),
    .B(_3691_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6874_ (.I(_1998_),
    .Z(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6875_ (.A1(_3798_),
    .A2(_1999_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6876_ (.A1(_1905_),
    .A2(_1994_),
    .A3(_2000_),
    .Z(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6877_ (.A1(_1979_),
    .A2(_1989_),
    .A3(_2001_),
    .Z(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6878_ (.A1(_1974_),
    .A2(_1976_),
    .A3(_2002_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6879_ (.A1(_1973_),
    .A2(_2003_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6880_ (.A1(_1970_),
    .A2(_2004_),
    .Z(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6881_ (.A1(_1956_),
    .A2(_1959_),
    .A3(_2005_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6882_ (.A1(_1939_),
    .A2(_1942_),
    .A3(_2006_),
    .Z(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6883_ (.A1(_1937_),
    .A2(_2007_),
    .ZN(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6884_ (.A1(_1934_),
    .A2(_2008_),
    .Z(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6885_ (.I(_2009_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6886_ (.I(\A[1][6] ),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6887_ (.A1(_2010_),
    .A2(_3776_),
    .A3(_1861_),
    .B1(_1698_),
    .B2(_3967_),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6888_ (.I(_2011_),
    .Z(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6889_ (.I(_2012_),
    .Z(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6890_ (.I(_2013_),
    .Z(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6891_ (.I(_2014_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6892_ (.A1(_1937_),
    .A2(_2007_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6893_ (.A1(_1934_),
    .A2(_2008_),
    .B(_2015_),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6894_ (.A1(_1942_),
    .A2(_2006_),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6895_ (.A1(_1942_),
    .A2(_2006_),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6896_ (.A1(_1939_),
    .A2(_2017_),
    .B(_2018_),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6897_ (.I(_1955_),
    .ZN(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6898_ (.A1(_1944_),
    .A2(_2020_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6899_ (.A1(_1945_),
    .A2(_1954_),
    .B(_2021_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6900_ (.A1(_1959_),
    .A2(_2005_),
    .Z(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6901_ (.A1(_1959_),
    .A2(_2005_),
    .Z(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6902_ (.A1(_1956_),
    .A2(_2023_),
    .B(_2024_),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6903_ (.A1(_4117_),
    .A2(_0012_),
    .A3(_1948_),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6904_ (.A1(_3510_),
    .A2(_0013_),
    .A3(_1951_),
    .ZN(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6905_ (.A1(_2026_),
    .A2(_2027_),
    .Z(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6906_ (.A1(_1960_),
    .A2(_1969_),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6907_ (.A1(_1965_),
    .A2(_1967_),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6908_ (.A1(_3776_),
    .A2(_3004_),
    .A3(_1754_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6909_ (.A1(_1878_),
    .A2(_2031_),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6910_ (.A1(_1966_),
    .A2(_2030_),
    .B(_2032_),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6911_ (.A1(_3903_),
    .A2(_1952_),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6912_ (.A1(_2033_),
    .A2(_2034_),
    .Z(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6913_ (.A1(_4227_),
    .A2(_2014_),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6914_ (.A1(_2035_),
    .A2(_2036_),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6915_ (.A1(_2029_),
    .A2(_2037_),
    .Z(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6916_ (.A1(_2028_),
    .A2(_2038_),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6917_ (.A1(_1973_),
    .A2(_2003_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6918_ (.A1(_1970_),
    .A2(_2004_),
    .B(_2040_),
    .ZN(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6919_ (.A1(_1964_),
    .A2(_1968_),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6920_ (.A1(_1974_),
    .A2(_1976_),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6921_ (.A1(_1961_),
    .A2(_1963_),
    .ZN(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6922_ (.I(_1862_),
    .Z(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6923_ (.A1(_4112_),
    .A2(_2045_),
    .ZN(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6924_ (.A1(_3792_),
    .A2(_2941_),
    .A3(_1807_),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6925_ (.A1(_2031_),
    .A2(_2047_),
    .Z(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6926_ (.A1(_2046_),
    .A2(_2048_),
    .Z(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6927_ (.I(_1744_),
    .Z(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6928_ (.A1(_3793_),
    .A2(_3861_),
    .A3(_2050_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6929_ (.A1(_4133_),
    .A2(_1882_),
    .ZN(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6930_ (.I(_4214_),
    .Z(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6931_ (.I(_1998_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6932_ (.I(_2054_),
    .Z(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6933_ (.A1(_2053_),
    .A2(_2055_),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6934_ (.A1(_2051_),
    .A2(_2052_),
    .A3(_2056_),
    .Z(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6935_ (.A1(_2044_),
    .A2(_2049_),
    .A3(_2057_),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6936_ (.A1(_2043_),
    .A2(_2058_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6937_ (.A1(_2042_),
    .A2(_2059_),
    .ZN(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6938_ (.A1(_1989_),
    .A2(_2001_),
    .Z(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6939_ (.A1(_1989_),
    .A2(_2001_),
    .ZN(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6940_ (.A1(_1974_),
    .A2(_1976_),
    .Z(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _6941_ (.A1(_1979_),
    .A2(_2061_),
    .A3(_2062_),
    .B1(_2002_),
    .B2(_2043_),
    .B3(_2063_),
    .ZN(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6942_ (.A1(_3969_),
    .A2(_1726_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6943_ (.A1(_3818_),
    .A2(_1907_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6944_ (.A1(_2065_),
    .A2(_2066_),
    .Z(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6945_ (.A1(_1984_),
    .A2(_2067_),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6946_ (.A1(_1991_),
    .A2(_1993_),
    .A3(_2000_),
    .Z(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6947_ (.A1(_1991_),
    .A2(_1993_),
    .B(_2000_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6948_ (.I(_1906_),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6949_ (.A1(_2069_),
    .A2(_2070_),
    .B(_2071_),
    .ZN(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6950_ (.A1(_1989_),
    .A2(_2001_),
    .B(_2072_),
    .ZN(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6951_ (.A1(_1985_),
    .A2(_1894_),
    .ZN(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6952_ (.A1(_2745_),
    .A2(_1777_),
    .B(\A[0][6] ),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6953_ (.A1(_3562_),
    .A2(_1848_),
    .ZN(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6954_ (.A1(_2075_),
    .A2(_2076_),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6955_ (.A1(_3832_),
    .A2(_2077_),
    .ZN(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6956_ (.A1(_4003_),
    .A2(_1770_),
    .B1(_1990_),
    .B2(_4088_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6957_ (.A1(_2079_),
    .A2(_2000_),
    .B(_1991_),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6958_ (.A1(_1178_),
    .A2(\C[1][6] ),
    .ZN(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6959_ (.A1(_3950_),
    .A2(_1971_),
    .A3(_2081_),
    .ZN(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6960_ (.A1(_3926_),
    .A2(_2081_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6961_ (.A1(_3998_),
    .A2(_1781_),
    .B(_2083_),
    .ZN(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6962_ (.A1(_2082_),
    .A2(_2084_),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6963_ (.A1(_1981_),
    .A2(_1982_),
    .B(_3990_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6964_ (.I(_2086_),
    .Z(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6965_ (.A1(_4157_),
    .A2(_2087_),
    .ZN(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6966_ (.A1(_2080_),
    .A2(_2085_),
    .A3(_2088_),
    .ZN(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6967_ (.A1(_2074_),
    .A2(_2078_),
    .A3(_2089_),
    .ZN(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6968_ (.A1(_2068_),
    .A2(_2073_),
    .A3(_2090_),
    .Z(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6969_ (.A1(_2064_),
    .A2(_2091_),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6970_ (.A1(_2060_),
    .A2(_2092_),
    .Z(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6971_ (.A1(_2039_),
    .A2(_2041_),
    .A3(_2093_),
    .Z(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6972_ (.A1(_2022_),
    .A2(_2025_),
    .A3(_2094_),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6973_ (.A1(_2016_),
    .A2(_2019_),
    .A3(_2095_),
    .Z(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6974_ (.I(_2096_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6975_ (.A1(net12),
    .A2(_1861_),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6976_ (.A1(\A[1][7] ),
    .A2(_3709_),
    .A3(_1743_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6977_ (.A1(_2097_),
    .A2(_2098_),
    .Z(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6978_ (.I(_2099_),
    .Z(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6979_ (.I(_2100_),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6980_ (.I(_2101_),
    .Z(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6981_ (.I(_2102_),
    .Z(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6982_ (.I(_2103_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6983_ (.A1(_2019_),
    .A2(_2095_),
    .ZN(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6984_ (.A1(_2019_),
    .A2(_2095_),
    .ZN(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6985_ (.A1(_2016_),
    .A2(_2104_),
    .B(_2105_),
    .ZN(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6986_ (.I(_2022_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6987_ (.A1(_2025_),
    .A2(_2094_),
    .Z(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6988_ (.A1(_2025_),
    .A2(_2094_),
    .Z(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6989_ (.A1(_2107_),
    .A2(_2108_),
    .B(_2109_),
    .ZN(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _6990_ (.A1(_1960_),
    .A2(_1969_),
    .A3(_2037_),
    .B1(_2038_),
    .B2(_2028_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6991_ (.A1(_2041_),
    .A2(_2093_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6992_ (.A1(_2041_),
    .A2(_2093_),
    .ZN(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6993_ (.A1(_2039_),
    .A2(_2112_),
    .B(_2113_),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6994_ (.A1(_0202_),
    .A2(_0013_),
    .A3(_2033_),
    .ZN(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6995_ (.A1(_2035_),
    .A2(_2036_),
    .B(_2115_),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6996_ (.A1(_2043_),
    .A2(_2058_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6997_ (.A1(_2042_),
    .A2(_2059_),
    .B(_2117_),
    .ZN(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6998_ (.A1(_2031_),
    .A2(_2047_),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6999_ (.I(_1949_),
    .Z(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7000_ (.A1(_4113_),
    .A2(_2120_),
    .A3(_2048_),
    .ZN(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7001_ (.A1(_2119_),
    .A2(_2121_),
    .ZN(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7002_ (.I(_2013_),
    .Z(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7003_ (.A1(_3229_),
    .A2(_2123_),
    .ZN(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7004_ (.A1(_2122_),
    .A2(_2124_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7005_ (.I(_2102_),
    .Z(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7006_ (.A1(_3888_),
    .A2(_2126_),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7007_ (.A1(_2125_),
    .A2(_2127_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7008_ (.A1(_2118_),
    .A2(_2128_),
    .Z(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7009_ (.A1(_2116_),
    .A2(_2129_),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7010_ (.A1(_2064_),
    .A2(_2091_),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7011_ (.A1(_2060_),
    .A2(_2092_),
    .B(_2131_),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7012_ (.A1(_2072_),
    .A2(_2061_),
    .A3(_2090_),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7013_ (.A1(_2072_),
    .A2(_2061_),
    .B(_2090_),
    .ZN(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7014_ (.A1(_2068_),
    .A2(_2133_),
    .B(_2134_),
    .ZN(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7015_ (.A1(_2065_),
    .A2(_2066_),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7016_ (.A1(_2074_),
    .A2(_2078_),
    .ZN(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7017_ (.A1(_4135_),
    .A2(_1882_),
    .ZN(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7018_ (.I(_2054_),
    .Z(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7019_ (.A1(_3816_),
    .A2(_2139_),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7020_ (.A1(_3980_),
    .A2(_1971_),
    .ZN(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7021_ (.A1(_2138_),
    .A2(_2140_),
    .A3(_2141_),
    .Z(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7022_ (.A1(_2137_),
    .A2(_2142_),
    .ZN(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7023_ (.A1(_2136_),
    .A2(_2143_),
    .ZN(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7024_ (.A1(_2074_),
    .A2(_2078_),
    .Z(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7025_ (.A1(_2085_),
    .A2(_2088_),
    .Z(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _7026_ (.A1(_2137_),
    .A2(_2145_),
    .A3(_2089_),
    .B1(_2146_),
    .B2(_2080_),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7027_ (.A1(_1529_),
    .A2(_1726_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7028_ (.A1(_1985_),
    .A2(_1907_),
    .ZN(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7029_ (.A1(_3854_),
    .A2(_1777_),
    .B(\A[0][7] ),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7030_ (.A1(_3894_),
    .A2(_1733_),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7031_ (.A1(_2150_),
    .A2(_2151_),
    .Z(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7032_ (.A1(_4150_),
    .A2(_2152_),
    .Z(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7033_ (.A1(_2148_),
    .A2(_2149_),
    .A3(_2153_),
    .Z(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7034_ (.I(\B[1][5] ),
    .Z(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7035_ (.I(_2155_),
    .Z(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7036_ (.A1(_1372_),
    .A2(\C[1][6] ),
    .A3(_2156_),
    .A4(_1826_),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7037_ (.A1(_2084_),
    .A2(_2088_),
    .B(_2157_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7038_ (.A1(_4089_),
    .A2(\C[1][7] ),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7039_ (.A1(_4003_),
    .A2(_1791_),
    .A3(_2159_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7040_ (.A1(_3925_),
    .A2(_2159_),
    .ZN(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7041_ (.A1(_1018_),
    .A2(_1840_),
    .B(_2161_),
    .ZN(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7042_ (.A1(_2075_),
    .A2(_2076_),
    .B(_3100_),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7043_ (.I(_2163_),
    .Z(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7044_ (.A1(_1838_),
    .A2(_2164_),
    .ZN(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _7045_ (.A1(_2160_),
    .A2(_2162_),
    .A3(_2165_),
    .Z(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7046_ (.A1(_2160_),
    .A2(_2162_),
    .B(_2165_),
    .ZN(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7047_ (.A1(_2166_),
    .A2(_2167_),
    .ZN(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7048_ (.A1(_2154_),
    .A2(_2158_),
    .A3(_2168_),
    .Z(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7049_ (.A1(_2144_),
    .A2(_2147_),
    .A3(_2169_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7050_ (.A1(_2044_),
    .A2(_2057_),
    .ZN(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7051_ (.A1(_2044_),
    .A2(_2057_),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7052_ (.A1(_2049_),
    .A2(_2171_),
    .B(_2172_),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7053_ (.A1(_1984_),
    .A2(_2067_),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7054_ (.A1(_3991_),
    .A2(_2993_),
    .A3(_1807_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7055_ (.A1(_2438_),
    .A2(_1927_),
    .Z(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7056_ (.A1(_2963_),
    .A2(_1863_),
    .Z(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7057_ (.A1(_2175_),
    .A2(_2176_),
    .A3(_2177_),
    .Z(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7058_ (.I(_3866_),
    .Z(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7059_ (.A1(_2179_),
    .A2(_1823_),
    .B1(_1998_),
    .B2(_3785_),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _7060_ (.A1(_3785_),
    .A2(_3866_),
    .A3(_1700_),
    .A4(_1998_),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7061_ (.A1(_2051_),
    .A2(_2180_),
    .B(_2181_),
    .ZN(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7062_ (.A1(_3960_),
    .A2(_3861_),
    .A3(_1755_),
    .ZN(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7063_ (.A1(_3821_),
    .A2(_3866_),
    .A3(_2050_),
    .ZN(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7064_ (.I(_2086_),
    .Z(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7065_ (.A1(_4214_),
    .A2(_2185_),
    .Z(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7066_ (.A1(_2183_),
    .A2(_2184_),
    .A3(_2186_),
    .Z(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7067_ (.A1(_2178_),
    .A2(_2182_),
    .A3(_2187_),
    .Z(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7068_ (.A1(_2174_),
    .A2(_2188_),
    .Z(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7069_ (.A1(_2173_),
    .A2(net40),
    .Z(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7070_ (.A1(_2135_),
    .A2(_2170_),
    .A3(_2190_),
    .Z(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7071_ (.A1(_2130_),
    .A2(_2132_),
    .A3(_2191_),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7072_ (.A1(_2114_),
    .A2(_2192_),
    .Z(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7073_ (.A1(_2111_),
    .A2(_2193_),
    .Z(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7074_ (.A1(_2106_),
    .A2(_2110_),
    .A3(_2194_),
    .ZN(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7075_ (.I(_2195_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7076_ (.A1(_2118_),
    .A2(_2128_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7077_ (.A1(_2116_),
    .A2(_2129_),
    .ZN(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7078_ (.A1(_2196_),
    .A2(_2197_),
    .ZN(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7079_ (.A1(_2132_),
    .A2(_2191_),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7080_ (.A1(_2132_),
    .A2(_2191_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7081_ (.A1(_2130_),
    .A2(_2199_),
    .B(_2200_),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7082_ (.A1(_4116_),
    .A2(_0014_),
    .A3(_2122_),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7083_ (.I(_2126_),
    .Z(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7084_ (.A1(_3889_),
    .A2(_2203_),
    .A3(_2125_),
    .ZN(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7085_ (.A1(_2202_),
    .A2(_2204_),
    .ZN(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7086_ (.A1(_2173_),
    .A2(_2189_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7087_ (.A1(_2174_),
    .A2(_2188_),
    .B(_2206_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7088_ (.A1(_0059_),
    .A2(_2120_),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7089_ (.A1(_2175_),
    .A2(_2177_),
    .Z(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7090_ (.A1(_2176_),
    .A2(_2209_),
    .ZN(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7091_ (.A1(_3004_),
    .A2(_1814_),
    .A3(_2208_),
    .B(_2210_),
    .ZN(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7092_ (.A1(_3240_),
    .A2(_2126_),
    .ZN(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7093_ (.A1(_2211_),
    .A2(_2212_),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7094_ (.A1(_2207_),
    .A2(_2213_),
    .Z(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7095_ (.A1(_2205_),
    .A2(_2214_),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7096_ (.A1(_2135_),
    .A2(_2170_),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7097_ (.I(_2190_),
    .ZN(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7098_ (.A1(_2135_),
    .A2(_2170_),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7099_ (.A1(_2216_),
    .A2(_2217_),
    .B(_2218_),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7100_ (.I(_2187_),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7101_ (.A1(_2182_),
    .A2(_2187_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7102_ (.A1(_2178_),
    .A2(_2221_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7103_ (.A1(_2182_),
    .A2(_2220_),
    .B(_2222_),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7104_ (.A1(_2137_),
    .A2(_2142_),
    .ZN(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7105_ (.A1(_2136_),
    .A2(_2143_),
    .B(_2224_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7106_ (.A1(_4112_),
    .A2(_2012_),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7107_ (.A1(_3015_),
    .A2(_1863_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7108_ (.A1(_2952_),
    .A2(_1927_),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7109_ (.A1(_2227_),
    .A2(_2228_),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7110_ (.A1(_2226_),
    .A2(_2229_),
    .Z(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7111_ (.A1(_2184_),
    .A2(_2186_),
    .Z(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7112_ (.A1(_2184_),
    .A2(_2186_),
    .Z(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7113_ (.A1(_2183_),
    .A2(_2231_),
    .B(_2232_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7114_ (.A1(_3861_),
    .A2(_1808_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7115_ (.I(_1753_),
    .Z(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7116_ (.I(_1754_),
    .Z(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7117_ (.A1(_2236_),
    .A2(_2179_),
    .A3(_2237_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7118_ (.A1(_4214_),
    .A2(_2164_),
    .ZN(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7119_ (.A1(_2238_),
    .A2(_2239_),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7120_ (.A1(_2235_),
    .A2(_2240_),
    .Z(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7121_ (.A1(_2230_),
    .A2(_2234_),
    .A3(_2241_),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7122_ (.A1(_2225_),
    .A2(_2242_),
    .Z(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7123_ (.A1(_2223_),
    .A2(_2243_),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7124_ (.A1(_2147_),
    .A2(_2169_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7125_ (.A1(_2147_),
    .A2(_2169_),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7126_ (.A1(_2144_),
    .A2(_2246_),
    .B(_2247_),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7127_ (.I(_2055_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7128_ (.A1(_4076_),
    .A2(_0004_),
    .B(_2141_),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7129_ (.I(_1899_),
    .Z(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7130_ (.A1(_0043_),
    .A2(_2250_),
    .A3(_2141_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7131_ (.A1(_2138_),
    .A2(_2249_),
    .B(_2251_),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7132_ (.A1(_2148_),
    .A2(_2149_),
    .Z(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7133_ (.A1(_2148_),
    .A2(_2149_),
    .Z(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7134_ (.A1(_2253_),
    .A2(_2153_),
    .B(_2255_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7135_ (.I(_2185_),
    .Z(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7136_ (.A1(_3817_),
    .A2(_2257_),
    .ZN(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7137_ (.A1(_3968_),
    .A2(_1841_),
    .ZN(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7138_ (.A1(_2258_),
    .A2(_2259_),
    .Z(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7139_ (.A1(_4035_),
    .A2(_1746_),
    .ZN(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7140_ (.A1(_2260_),
    .A2(_2261_),
    .Z(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7141_ (.A1(_2256_),
    .A2(_2262_),
    .Z(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7142_ (.A1(_2252_),
    .A2(_2263_),
    .ZN(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7143_ (.A1(_2166_),
    .A2(_2167_),
    .B(_2158_),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7144_ (.A1(_2158_),
    .A2(_2166_),
    .A3(_2167_),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7145_ (.A1(_2154_),
    .A2(_2266_),
    .B(_2267_),
    .ZN(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _7146_ (.A1(_4001_),
    .A2(_1319_),
    .A3(_1980_),
    .A4(_1999_),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7147_ (.I(_2269_),
    .Z(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7148_ (.A1(_1530_),
    .A2(_1826_),
    .B1(_0004_),
    .B2(_4069_),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7149_ (.A1(_2270_),
    .A2(_2271_),
    .ZN(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7150_ (.A1(_4090_),
    .A2(\C[1][7] ),
    .A3(_2156_),
    .A4(_1840_),
    .ZN(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7151_ (.A1(_2162_),
    .A2(_2165_),
    .B(_2273_),
    .ZN(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7152_ (.I(_1902_),
    .Z(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7153_ (.A1(_3982_),
    .A2(\C[1][8] ),
    .A3(_2155_),
    .A4(_2275_),
    .Z(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7154_ (.A1(_0513_),
    .A2(\C[1][8] ),
    .A3(_2652_),
    .Z(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7155_ (.A1(_1018_),
    .A2(_2275_),
    .B(_2278_),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7156_ (.A1(_2277_),
    .A2(_2279_),
    .ZN(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7157_ (.A1(_2150_),
    .A2(_2151_),
    .B(_3991_),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7158_ (.I(_2281_),
    .Z(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7159_ (.A1(_1838_),
    .A2(_2282_),
    .ZN(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7160_ (.A1(_2274_),
    .A2(_2280_),
    .A3(_2283_),
    .Z(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7161_ (.A1(_2272_),
    .A2(_2284_),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7162_ (.A1(_2264_),
    .A2(_2268_),
    .A3(_2285_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7163_ (.A1(_2245_),
    .A2(_2248_),
    .A3(_2286_),
    .ZN(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7164_ (.A1(_2215_),
    .A2(_2219_),
    .A3(_2288_),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7165_ (.A1(_2201_),
    .A2(_2289_),
    .Z(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7166_ (.A1(_2198_),
    .A2(_2290_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7167_ (.A1(_2114_),
    .A2(_2192_),
    .Z(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7168_ (.A1(_2111_),
    .A2(_2193_),
    .B(_2292_),
    .ZN(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7169_ (.A1(_2291_),
    .A2(_2293_),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7170_ (.A1(_2110_),
    .A2(_2194_),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7171_ (.A1(_2016_),
    .A2(_2104_),
    .B1(_2110_),
    .B2(_2194_),
    .C(_2105_),
    .ZN(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7172_ (.A1(_2295_),
    .A2(_2296_),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7173_ (.A1(_2294_),
    .A2(_2297_),
    .ZN(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7174_ (.I(_2299_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7175_ (.A1(_2201_),
    .A2(_2289_),
    .Z(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7176_ (.A1(_2198_),
    .A2(_2290_),
    .B(_2300_),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7177_ (.A1(_2207_),
    .A2(_2213_),
    .ZN(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7178_ (.A1(_2205_),
    .A2(_2214_),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7179_ (.A1(_2302_),
    .A2(_2303_),
    .ZN(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7180_ (.A1(_2219_),
    .A2(_2288_),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7181_ (.A1(_2219_),
    .A2(_2288_),
    .ZN(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7182_ (.A1(_2215_),
    .A2(_2305_),
    .B(_2306_),
    .ZN(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7183_ (.A1(_0220_),
    .A2(_0015_),
    .A3(_2211_),
    .Z(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7184_ (.A1(_2225_),
    .A2(_2242_),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7185_ (.A1(_2223_),
    .A2(_2243_),
    .ZN(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7186_ (.A1(_2310_),
    .A2(_2311_),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7187_ (.A1(_3026_),
    .A2(_1929_),
    .ZN(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _7188_ (.A1(_2208_),
    .A2(_2313_),
    .B1(_2229_),
    .B2(_2226_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7189_ (.A1(_2312_),
    .A2(_2314_),
    .Z(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7190_ (.A1(_2309_),
    .A2(_2315_),
    .Z(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7191_ (.A1(_2248_),
    .A2(_2286_),
    .ZN(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7192_ (.A1(_2248_),
    .A2(_2286_),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7193_ (.A1(_2245_),
    .A2(_2317_),
    .B(_2318_),
    .ZN(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7194_ (.I(_2234_),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7195_ (.A1(_2321_),
    .A2(_2241_),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7196_ (.A1(_2234_),
    .A2(_2241_),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7197_ (.A1(_2230_),
    .A2(_2323_),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7198_ (.A1(_2322_),
    .A2(_2324_),
    .ZN(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7199_ (.A1(_2256_),
    .A2(_2262_),
    .Z(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7200_ (.A1(_2252_),
    .A2(_2263_),
    .B(_2326_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7201_ (.A1(_1768_),
    .A2(_2100_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7202_ (.A1(_4195_),
    .A2(_2012_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7203_ (.A1(_2313_),
    .A2(_2329_),
    .ZN(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7204_ (.A1(_2328_),
    .A2(_2331_),
    .Z(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7205_ (.A1(_2179_),
    .A2(_1757_),
    .A3(_2239_),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7206_ (.A1(_2235_),
    .A2(_2240_),
    .B(_2333_),
    .ZN(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7207_ (.A1(_3863_),
    .A2(_2045_),
    .ZN(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7208_ (.A1(_4133_),
    .A2(_1809_),
    .ZN(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7209_ (.A1(_2053_),
    .A2(_2282_),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7210_ (.A1(_2335_),
    .A2(_2336_),
    .A3(_2337_),
    .Z(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7211_ (.A1(_2334_),
    .A2(_2338_),
    .ZN(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7212_ (.A1(_2332_),
    .A2(_2339_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7213_ (.A1(_2327_),
    .A2(_2340_),
    .Z(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7214_ (.A1(_2325_),
    .A2(_2342_),
    .Z(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7215_ (.A1(_2268_),
    .A2(_2285_),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7216_ (.A1(_2268_),
    .A2(_2285_),
    .ZN(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7217_ (.A1(_2264_),
    .A2(_2344_),
    .B(_2345_),
    .ZN(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7218_ (.A1(_2258_),
    .A2(_2259_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7219_ (.A1(_2260_),
    .A2(_2261_),
    .B(_2347_),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7220_ (.A1(_4035_),
    .A2(_1757_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7221_ (.I(_2164_),
    .Z(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7222_ (.A1(_3817_),
    .A2(_2350_),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7223_ (.I(_1962_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7224_ (.A1(_3969_),
    .A2(_0003_),
    .ZN(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7225_ (.A1(_2349_),
    .A2(_2351_),
    .A3(_2353_),
    .Z(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7226_ (.A1(_2270_),
    .A2(_2348_),
    .A3(_2354_),
    .Z(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7227_ (.A1(_2280_),
    .A2(_2283_),
    .Z(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7228_ (.I(_2274_),
    .ZN(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7229_ (.A1(_2269_),
    .A2(_2271_),
    .A3(_2284_),
    .B1(_2356_),
    .B2(_2357_),
    .ZN(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7230_ (.A1(_1985_),
    .A2(_1529_),
    .A3(_1975_),
    .A4(_2087_),
    .ZN(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7231_ (.A1(_1319_),
    .A2(_1791_),
    .B1(_1983_),
    .B2(_1163_),
    .ZN(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7232_ (.A1(_2359_),
    .A2(_2360_),
    .ZN(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7233_ (.A1(_0514_),
    .A2(\C[1][8] ),
    .A3(_2156_),
    .A4(_1903_),
    .ZN(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7234_ (.A1(_2279_),
    .A2(_2283_),
    .B(_2363_),
    .ZN(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7235_ (.A1(_3957_),
    .A2(_2139_),
    .ZN(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7236_ (.A1(_4090_),
    .A2(\C[1][9] ),
    .A3(_3974_),
    .ZN(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7237_ (.A1(_1178_),
    .A2(\C[1][9] ),
    .A3(_2155_),
    .A4(_2139_),
    .Z(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7238_ (.A1(_2365_),
    .A2(_2366_),
    .B(_2367_),
    .ZN(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7239_ (.A1(_2364_),
    .A2(_2368_),
    .ZN(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7240_ (.A1(_2361_),
    .A2(_2369_),
    .Z(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7241_ (.A1(_2358_),
    .A2(_2370_),
    .ZN(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7242_ (.A1(_2355_),
    .A2(_2371_),
    .Z(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7243_ (.A1(_2346_),
    .A2(_2372_),
    .Z(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7244_ (.A1(_2343_),
    .A2(_2374_),
    .Z(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7245_ (.A1(_2320_),
    .A2(_2375_),
    .Z(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7246_ (.A1(_2316_),
    .A2(_2376_),
    .Z(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7247_ (.A1(_2304_),
    .A2(_2307_),
    .A3(_2377_),
    .ZN(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7248_ (.A1(_2301_),
    .A2(_2378_),
    .ZN(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7249_ (.A1(_2295_),
    .A2(_2294_),
    .A3(_2296_),
    .B1(_2291_),
    .B2(_2293_),
    .ZN(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7250_ (.A1(_2379_),
    .A2(_2380_),
    .ZN(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7251_ (.I(_2381_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7252_ (.A1(_2312_),
    .A2(_2314_),
    .ZN(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7253_ (.A1(_2309_),
    .A2(_2315_),
    .ZN(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7254_ (.A1(_2382_),
    .A2(_2384_),
    .ZN(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7255_ (.A1(_2320_),
    .A2(_2375_),
    .Z(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7256_ (.A1(_2316_),
    .A2(_2376_),
    .B(_2386_),
    .ZN(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7257_ (.A1(_2325_),
    .A2(_2342_),
    .ZN(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7258_ (.A1(_2327_),
    .A2(_2340_),
    .B(_2388_),
    .ZN(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7259_ (.I(_2100_),
    .Z(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7260_ (.A1(_1768_),
    .A2(_2390_),
    .A3(_2331_),
    .B1(_2329_),
    .B2(_2313_),
    .ZN(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7261_ (.A1(_2389_),
    .A2(_2391_),
    .ZN(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7262_ (.A1(_2346_),
    .A2(_2372_),
    .Z(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7263_ (.A1(_2343_),
    .A2(_2374_),
    .B(_2393_),
    .ZN(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7264_ (.A1(_2334_),
    .A2(_2338_),
    .Z(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7265_ (.A1(_2332_),
    .A2(_2339_),
    .B(_2396_),
    .ZN(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7266_ (.A1(_2270_),
    .A2(_2354_),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7267_ (.A1(_2270_),
    .A2(_2354_),
    .ZN(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7268_ (.A1(_2348_),
    .A2(_2398_),
    .B(_2399_),
    .ZN(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7269_ (.A1(_4133_),
    .A2(_1864_),
    .ZN(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7270_ (.A1(_3864_),
    .A2(_1928_),
    .ZN(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7271_ (.A1(_2401_),
    .A2(_2402_),
    .Z(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7272_ (.I(_2282_),
    .Z(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7273_ (.A1(_3873_),
    .A2(_1810_),
    .B1(_2404_),
    .B2(_2053_),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7274_ (.A1(_2053_),
    .A2(_3873_),
    .A3(_1810_),
    .A4(_2404_),
    .ZN(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7275_ (.A1(_2335_),
    .A2(_2406_),
    .B(_2407_),
    .ZN(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7276_ (.A1(_2403_),
    .A2(_2408_),
    .Z(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7277_ (.A1(_0980_),
    .A2(_2101_),
    .ZN(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7278_ (.A1(_2329_),
    .A2(_2410_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7279_ (.A1(_0060_),
    .A2(_2013_),
    .B1(_2102_),
    .B2(_0059_),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7280_ (.A1(_2411_),
    .A2(_2412_),
    .ZN(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7281_ (.A1(_2409_),
    .A2(_2413_),
    .Z(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7282_ (.A1(_2400_),
    .A2(_2414_),
    .Z(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7283_ (.A1(_2397_),
    .A2(_2415_),
    .ZN(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7284_ (.A1(_2358_),
    .A2(_2370_),
    .ZN(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7285_ (.A1(_2355_),
    .A2(_2371_),
    .B(_2418_),
    .ZN(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7286_ (.A1(_2351_),
    .A2(_2353_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7287_ (.A1(_2351_),
    .A2(_2353_),
    .ZN(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7288_ (.A1(_2349_),
    .A2(_2420_),
    .B(_2421_),
    .ZN(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7289_ (.A1(_4034_),
    .A2(_1808_),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7290_ (.A1(_3816_),
    .A2(_2281_),
    .ZN(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7291_ (.A1(_3968_),
    .A2(_2139_),
    .ZN(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7292_ (.A1(_2424_),
    .A2(_2425_),
    .Z(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7293_ (.A1(_2423_),
    .A2(_2426_),
    .Z(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7294_ (.A1(_2359_),
    .A2(_2428_),
    .Z(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7295_ (.A1(_2422_),
    .A2(_2429_),
    .Z(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7296_ (.A1(_2364_),
    .A2(_2368_),
    .ZN(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7297_ (.A1(_2364_),
    .A2(_2368_),
    .ZN(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7298_ (.A1(_2361_),
    .A2(_2431_),
    .B(_2432_),
    .ZN(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7299_ (.A1(_1018_),
    .A2(_2257_),
    .ZN(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7300_ (.A1(_0473_),
    .A2(\C[1][10] ),
    .A3(_3974_),
    .ZN(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7301_ (.A1(_3971_),
    .A2(\C[1][10] ),
    .A3(_2155_),
    .A4(_2185_),
    .Z(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7302_ (.A1(_2434_),
    .A2(_2435_),
    .B(_2436_),
    .ZN(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7303_ (.A1(_2367_),
    .A2(_2437_),
    .Z(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7304_ (.A1(_3917_),
    .A2(_2350_),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7305_ (.A1(_4085_),
    .A2(_1962_),
    .ZN(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7306_ (.A1(_2440_),
    .A2(_2441_),
    .Z(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7307_ (.A1(_2439_),
    .A2(_2442_),
    .Z(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7308_ (.A1(_2433_),
    .A2(_2443_),
    .Z(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7309_ (.A1(_2430_),
    .A2(_2444_),
    .Z(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7310_ (.A1(_2419_),
    .A2(_2445_),
    .ZN(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7311_ (.A1(_2417_),
    .A2(_2446_),
    .ZN(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7312_ (.A1(_2395_),
    .A2(_2447_),
    .ZN(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7313_ (.A1(_2392_),
    .A2(_2448_),
    .ZN(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7314_ (.A1(_2387_),
    .A2(_2450_),
    .Z(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7315_ (.A1(_2385_),
    .A2(_2451_),
    .ZN(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7316_ (.A1(_2307_),
    .A2(_2377_),
    .Z(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7317_ (.A1(_2307_),
    .A2(_2377_),
    .Z(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7318_ (.A1(_2304_),
    .A2(_2453_),
    .B(_2454_),
    .ZN(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7319_ (.A1(_2452_),
    .A2(_2455_),
    .Z(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _7320_ (.A1(_2295_),
    .A2(_2294_),
    .A3(_2296_),
    .A4(_2379_),
    .Z(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7321_ (.A1(_2291_),
    .A2(_2293_),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7322_ (.A1(_2301_),
    .A2(_2378_),
    .ZN(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7323_ (.A1(_2301_),
    .A2(_2378_),
    .ZN(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7324_ (.A1(_2458_),
    .A2(_2459_),
    .B(_2461_),
    .ZN(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7325_ (.A1(_2457_),
    .A2(_2462_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7326_ (.A1(_2456_),
    .A2(_2463_),
    .Z(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7327_ (.I(_2464_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7328_ (.A1(_2387_),
    .A2(_2450_),
    .ZN(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7329_ (.A1(_2385_),
    .A2(_2451_),
    .B(_2465_),
    .ZN(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7330_ (.A1(_2389_),
    .A2(_2391_),
    .ZN(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7331_ (.A1(_2395_),
    .A2(_2447_),
    .Z(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7332_ (.A1(_2392_),
    .A2(_2448_),
    .B(_2468_),
    .ZN(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7333_ (.A1(_2400_),
    .A2(_2414_),
    .ZN(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7334_ (.A1(_2397_),
    .A2(_2415_),
    .ZN(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7335_ (.A1(_2471_),
    .A2(_2472_),
    .ZN(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7336_ (.A1(_2411_),
    .A2(_2473_),
    .Z(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7337_ (.A1(_2419_),
    .A2(_2445_),
    .ZN(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7338_ (.A1(_2417_),
    .A2(_2446_),
    .B(_2475_),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7339_ (.A1(_2403_),
    .A2(_2408_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7340_ (.A1(_2409_),
    .A2(_2413_),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7341_ (.A1(_2477_),
    .A2(_2478_),
    .ZN(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7342_ (.I(_2359_),
    .ZN(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7343_ (.A1(_2480_),
    .A2(_2428_),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7344_ (.A1(_2422_),
    .A2(_2429_),
    .B(_2482_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7345_ (.A1(_3877_),
    .A2(_2123_),
    .ZN(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7346_ (.A1(_3874_),
    .A2(_1952_),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7347_ (.A1(_3877_),
    .A2(_2120_),
    .B(_2485_),
    .ZN(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7348_ (.A1(_2484_),
    .A2(_2486_),
    .Z(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7349_ (.A1(_2410_),
    .A2(_2487_),
    .Z(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7350_ (.A1(_2483_),
    .A2(_2488_),
    .Z(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7351_ (.A1(_2479_),
    .A2(_2489_),
    .Z(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7352_ (.A1(_2433_),
    .A2(_2443_),
    .Z(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7353_ (.A1(_2430_),
    .A2(_2444_),
    .B(_2491_),
    .ZN(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7354_ (.A1(_2367_),
    .A2(_2437_),
    .Z(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7355_ (.A1(_2439_),
    .A2(_2442_),
    .B(_2494_),
    .ZN(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7356_ (.A1(_3998_),
    .A2(_2350_),
    .ZN(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7357_ (.A1(_1247_),
    .A2(\C[1][11] ),
    .A3(_0476_),
    .ZN(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7358_ (.A1(_4090_),
    .A2(\C[1][11] ),
    .A3(_2156_),
    .A4(_2164_),
    .Z(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7359_ (.A1(_2496_),
    .A2(_2497_),
    .B(_2498_),
    .ZN(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7360_ (.A1(_2436_),
    .A2(_2499_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7361_ (.I(_2282_),
    .Z(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7362_ (.A1(_4069_),
    .A2(_1529_),
    .A3(_0004_),
    .A4(_2501_),
    .ZN(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7363_ (.A1(_1319_),
    .A2(_1999_),
    .B1(_2152_),
    .B2(_1164_),
    .ZN(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7364_ (.A1(_2502_),
    .A2(_2504_),
    .ZN(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7365_ (.A1(_2500_),
    .A2(_2505_),
    .ZN(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7366_ (.A1(_2495_),
    .A2(_2506_),
    .ZN(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7367_ (.A1(_2424_),
    .A2(_2425_),
    .ZN(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7368_ (.A1(_2423_),
    .A2(_2426_),
    .B(_2508_),
    .ZN(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7369_ (.A1(_2440_),
    .A2(_2441_),
    .Z(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7370_ (.A1(_1295_),
    .A2(_1949_),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7371_ (.I(_2087_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7372_ (.A1(_1538_),
    .A2(_0005_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7373_ (.A1(_2510_),
    .A2(_2511_),
    .A3(_2512_),
    .Z(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7374_ (.A1(_2509_),
    .A2(_2514_),
    .ZN(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7375_ (.A1(_2507_),
    .A2(_2515_),
    .ZN(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7376_ (.A1(_2493_),
    .A2(_2516_),
    .Z(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7377_ (.A1(_2490_),
    .A2(_2517_),
    .Z(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7378_ (.A1(_2476_),
    .A2(_2518_),
    .Z(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7379_ (.A1(_2474_),
    .A2(_2519_),
    .Z(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7380_ (.A1(_2467_),
    .A2(_2469_),
    .A3(_2520_),
    .ZN(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7381_ (.A1(_2466_),
    .A2(_2521_),
    .Z(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7382_ (.A1(_2452_),
    .A2(_2455_),
    .Z(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7383_ (.A1(_2456_),
    .A2(_2463_),
    .ZN(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7384_ (.A1(_2523_),
    .A2(_2525_),
    .ZN(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7385_ (.A1(_2522_),
    .A2(_2526_),
    .ZN(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7386_ (.I(_2527_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7387_ (.A1(_2452_),
    .A2(_2455_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7388_ (.A1(_2457_),
    .A2(_2462_),
    .B(_2522_),
    .C(_2528_),
    .ZN(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7389_ (.A1(_2385_),
    .A2(_2451_),
    .Z(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7390_ (.A1(_2465_),
    .A2(_2530_),
    .A3(_2521_),
    .ZN(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7391_ (.A1(_2465_),
    .A2(_2530_),
    .B(_2521_),
    .ZN(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7392_ (.A1(_2523_),
    .A2(_2531_),
    .B(_2532_),
    .ZN(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7393_ (.A1(_2529_),
    .A2(_2533_),
    .ZN(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7394_ (.A1(_2411_),
    .A2(_2473_),
    .Z(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7395_ (.A1(_2476_),
    .A2(_2518_),
    .ZN(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7396_ (.A1(_2474_),
    .A2(_2519_),
    .ZN(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7397_ (.A1(_2537_),
    .A2(_2538_),
    .ZN(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7398_ (.A1(_2483_),
    .A2(_2488_),
    .ZN(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7399_ (.A1(_2479_),
    .A2(_2489_),
    .ZN(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7400_ (.A1(_2540_),
    .A2(_2541_),
    .ZN(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7401_ (.A1(_2490_),
    .A2(_2517_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7402_ (.A1(_2493_),
    .A2(_2516_),
    .B(_2543_),
    .ZN(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7403_ (.A1(_2495_),
    .A2(_2506_),
    .ZN(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7404_ (.A1(_2507_),
    .A2(_2515_),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7405_ (.A1(_2546_),
    .A2(_2547_),
    .ZN(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7406_ (.A1(_2500_),
    .A2(_2505_),
    .ZN(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7407_ (.A1(_2436_),
    .A2(_2499_),
    .B(_2549_),
    .ZN(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7408_ (.A1(_1530_),
    .A2(_0005_),
    .ZN(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7409_ (.A1(_3999_),
    .A2(_2404_),
    .Z(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7410_ (.A1(\C[1][12] ),
    .A2(_3929_),
    .Z(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7411_ (.A1(_1372_),
    .A2(\C[1][12] ),
    .A3(_2552_),
    .ZN(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7412_ (.A1(_2552_),
    .A2(_2553_),
    .B(_2554_),
    .ZN(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7413_ (.A1(_2498_),
    .A2(_2555_),
    .Z(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7414_ (.A1(_2550_),
    .A2(_2551_),
    .A3(_2557_),
    .Z(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7415_ (.A1(_2511_),
    .A2(_2512_),
    .Z(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7416_ (.I(_2502_),
    .ZN(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7417_ (.A1(_1295_),
    .A2(_1930_),
    .ZN(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7418_ (.I(_2163_),
    .Z(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7419_ (.A1(_1538_),
    .A2(_2562_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7420_ (.A1(_2561_),
    .A2(_2563_),
    .Z(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7421_ (.A1(_2560_),
    .A2(_2564_),
    .Z(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7422_ (.A1(_2559_),
    .A2(_2565_),
    .Z(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7423_ (.A1(_2558_),
    .A2(_2566_),
    .ZN(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7424_ (.A1(_2548_),
    .A2(_2568_),
    .Z(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7425_ (.A1(_0061_),
    .A2(_2014_),
    .Z(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7426_ (.A1(_2335_),
    .A2(_2485_),
    .A3(_2570_),
    .ZN(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7427_ (.A1(_2410_),
    .A2(_2487_),
    .ZN(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7428_ (.A1(_2571_),
    .A2(_2572_),
    .ZN(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7429_ (.I(_2559_),
    .ZN(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7430_ (.A1(_2511_),
    .A2(_2512_),
    .Z(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7431_ (.A1(_2510_),
    .A2(_2574_),
    .A3(_2575_),
    .B1(_2514_),
    .B2(_2509_),
    .ZN(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7432_ (.A1(_3883_),
    .A2(_2126_),
    .ZN(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7433_ (.I(_2123_),
    .Z(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7434_ (.A1(_0062_),
    .A2(_2579_),
    .A3(_2402_),
    .ZN(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7435_ (.A1(_2577_),
    .A2(_2580_),
    .Z(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7436_ (.A1(_2576_),
    .A2(_2581_),
    .ZN(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7437_ (.A1(_2573_),
    .A2(_2582_),
    .Z(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7438_ (.A1(_2569_),
    .A2(_2583_),
    .Z(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7439_ (.A1(_2544_),
    .A2(_2584_),
    .Z(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7440_ (.A1(_2542_),
    .A2(_2585_),
    .Z(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7441_ (.A1(_2539_),
    .A2(_2586_),
    .Z(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7442_ (.A1(_2536_),
    .A2(_2587_),
    .Z(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7443_ (.A1(_2469_),
    .A2(_2520_),
    .ZN(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7444_ (.A1(_2469_),
    .A2(_2520_),
    .ZN(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7445_ (.A1(_2467_),
    .A2(_2590_),
    .B(_2591_),
    .ZN(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7446_ (.A1(_2588_),
    .A2(_2592_),
    .Z(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7447_ (.A1(_2535_),
    .A2(_2593_),
    .ZN(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7448_ (.I(_2594_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7449_ (.A1(_2576_),
    .A2(_2581_),
    .ZN(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7450_ (.A1(_2573_),
    .A2(_2582_),
    .B(_2595_),
    .ZN(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7451_ (.A1(_2548_),
    .A2(_2568_),
    .ZN(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7452_ (.A1(_2569_),
    .A2(_2583_),
    .B(_2597_),
    .ZN(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7453_ (.A1(_2560_),
    .A2(_2564_),
    .ZN(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7454_ (.A1(_2574_),
    .A2(_2565_),
    .ZN(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7455_ (.A1(_2600_),
    .A2(_2601_),
    .ZN(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7456_ (.A1(_2485_),
    .A2(_2484_),
    .ZN(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7457_ (.A1(_2179_),
    .A2(_2390_),
    .ZN(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7458_ (.A1(_2103_),
    .A2(_2570_),
    .ZN(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7459_ (.A1(_2603_),
    .A2(_2604_),
    .B(_2605_),
    .ZN(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7460_ (.A1(_2602_),
    .A2(_2606_),
    .ZN(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7461_ (.A1(_2551_),
    .A2(_2557_),
    .ZN(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7462_ (.A1(_2551_),
    .A2(_2557_),
    .Z(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7463_ (.A1(_2550_),
    .A2(_2608_),
    .A3(_2609_),
    .B1(_2558_),
    .B2(_2566_),
    .ZN(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7464_ (.A1(_2561_),
    .A2(_2563_),
    .ZN(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7465_ (.A1(_1419_),
    .A2(_2579_),
    .ZN(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7466_ (.I(_2501_),
    .Z(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7467_ (.A1(_1538_),
    .A2(_2614_),
    .ZN(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7468_ (.A1(_2613_),
    .A2(_2615_),
    .Z(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7469_ (.A1(_2613_),
    .A2(_2615_),
    .Z(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7470_ (.I(_2617_),
    .ZN(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7471_ (.A1(_2616_),
    .A2(_2618_),
    .ZN(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7472_ (.A1(_2612_),
    .A2(_2619_),
    .ZN(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7473_ (.I(_2498_),
    .ZN(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7474_ (.A1(_1533_),
    .A2(_1983_),
    .A3(_2557_),
    .B1(_2555_),
    .B2(_2622_),
    .ZN(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7475_ (.A1(\C[1][13] ),
    .A2(_0185_),
    .ZN(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7476_ (.A1(_2554_),
    .A2(_2624_),
    .ZN(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7477_ (.A1(\C[1][12] ),
    .A2(\C[1][13] ),
    .A3(_0185_),
    .A4(_2552_),
    .ZN(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7478_ (.A1(_2625_),
    .A2(_2626_),
    .ZN(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7479_ (.I(_2562_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7480_ (.A1(_1530_),
    .A2(_0006_),
    .Z(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7481_ (.A1(_2627_),
    .A2(_2628_),
    .ZN(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7482_ (.A1(_2623_),
    .A2(_2629_),
    .Z(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7483_ (.A1(_2620_),
    .A2(_2630_),
    .Z(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7484_ (.A1(_2611_),
    .A2(_2632_),
    .ZN(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7485_ (.A1(_2607_),
    .A2(_2633_),
    .Z(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7486_ (.A1(_2598_),
    .A2(_2634_),
    .Z(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7487_ (.A1(_2596_),
    .A2(_2635_),
    .ZN(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7488_ (.A1(_2544_),
    .A2(_2584_),
    .ZN(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7489_ (.A1(_2542_),
    .A2(_2585_),
    .ZN(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7490_ (.A1(_2637_),
    .A2(_2638_),
    .ZN(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7491_ (.A1(_2636_),
    .A2(_2639_),
    .Z(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7492_ (.A1(_2539_),
    .A2(_2586_),
    .ZN(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7493_ (.A1(_2536_),
    .A2(_2587_),
    .ZN(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7494_ (.A1(_2641_),
    .A2(_2643_),
    .ZN(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7495_ (.A1(_2588_),
    .A2(_2592_),
    .ZN(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7496_ (.A1(_2529_),
    .A2(_2533_),
    .B(_2593_),
    .ZN(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7497_ (.A1(_2645_),
    .A2(_2646_),
    .ZN(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7498_ (.A1(_2640_),
    .A2(_2644_),
    .A3(_2647_),
    .ZN(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7499_ (.I(_2648_),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7500_ (.I(_2636_),
    .ZN(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7501_ (.A1(_2649_),
    .A2(_2639_),
    .ZN(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7502_ (.A1(_2603_),
    .A2(_2604_),
    .B(_2605_),
    .C(_2602_),
    .ZN(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7503_ (.I(_2607_),
    .ZN(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7504_ (.A1(_2611_),
    .A2(_2632_),
    .ZN(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7505_ (.A1(_2653_),
    .A2(_2633_),
    .B(_2654_),
    .ZN(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7506_ (.A1(_2623_),
    .A2(_2629_),
    .ZN(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7507_ (.A1(_2620_),
    .A2(_2630_),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7508_ (.A1(_2656_),
    .A2(_2657_),
    .ZN(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7509_ (.A1(_2100_),
    .A2(_2616_),
    .Z(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7510_ (.A1(_4035_),
    .A2(_2390_),
    .B(_2616_),
    .ZN(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7511_ (.A1(_2659_),
    .A2(_2660_),
    .ZN(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7512_ (.A1(_2625_),
    .A2(_2626_),
    .A3(_2628_),
    .ZN(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7513_ (.A1(_2626_),
    .A2(_2662_),
    .Z(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7514_ (.I(_2501_),
    .Z(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7515_ (.A1(_1597_),
    .A2(\C[1][14] ),
    .A3(\B[1][7] ),
    .A4(_2665_),
    .ZN(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7516_ (.A1(\C[1][14] ),
    .A2(_0186_),
    .ZN(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7517_ (.A1(_1533_),
    .A2(_2152_),
    .B(_2667_),
    .ZN(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7518_ (.A1(_2666_),
    .A2(_2668_),
    .ZN(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7519_ (.A1(_2664_),
    .A2(_2669_),
    .ZN(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7520_ (.A1(_2661_),
    .A2(_2670_),
    .Z(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7521_ (.A1(_2658_),
    .A2(_2671_),
    .Z(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7522_ (.A1(_2612_),
    .A2(_2616_),
    .A3(_2618_),
    .ZN(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7523_ (.A1(_2570_),
    .A2(_2604_),
    .ZN(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7524_ (.A1(_2673_),
    .A2(_2675_),
    .Z(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7525_ (.A1(_2672_),
    .A2(_2676_),
    .Z(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7526_ (.A1(_2651_),
    .A2(_2655_),
    .A3(_2677_),
    .ZN(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7527_ (.A1(_2598_),
    .A2(_2634_),
    .ZN(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7528_ (.A1(_2596_),
    .A2(_2635_),
    .B(_2679_),
    .ZN(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7529_ (.A1(_2678_),
    .A2(_2680_),
    .Z(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7530_ (.A1(_2650_),
    .A2(_2681_),
    .Z(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7531_ (.A1(_2641_),
    .A2(_2643_),
    .B(_2640_),
    .ZN(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7532_ (.A1(_2588_),
    .A2(_2592_),
    .B(_2683_),
    .ZN(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7533_ (.A1(_2641_),
    .A2(_2643_),
    .A3(_2640_),
    .ZN(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7534_ (.I(_2686_),
    .ZN(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7535_ (.A1(_2646_),
    .A2(_2684_),
    .B(_2687_),
    .ZN(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7536_ (.A1(_2682_),
    .A2(_2688_),
    .Z(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7537_ (.I(_2689_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7538_ (.A1(_2650_),
    .A2(_2681_),
    .ZN(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7539_ (.A1(_2682_),
    .A2(_2688_),
    .B(_2690_),
    .ZN(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7540_ (.I(_2680_),
    .ZN(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7541_ (.A1(_2678_),
    .A2(_2692_),
    .ZN(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7542_ (.A1(_2673_),
    .A2(_2675_),
    .ZN(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7543_ (.A1(_2655_),
    .A2(_2677_),
    .ZN(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7544_ (.A1(_2655_),
    .A2(_2677_),
    .ZN(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7545_ (.A1(_2651_),
    .A2(_2696_),
    .B(_2697_),
    .ZN(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7546_ (.A1(_2658_),
    .A2(_2671_),
    .ZN(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7547_ (.A1(_2672_),
    .A2(_2676_),
    .ZN(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7548_ (.A1(_2699_),
    .A2(_2700_),
    .ZN(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7549_ (.A1(_2664_),
    .A2(_2669_),
    .ZN(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7550_ (.A1(_2661_),
    .A2(_2670_),
    .ZN(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7551_ (.A1(\C[1][15] ),
    .A2(_0947_),
    .ZN(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7552_ (.A1(\C[1][15] ),
    .A2(_1630_),
    .ZN(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7553_ (.A1(_2666_),
    .A2(_2705_),
    .ZN(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7554_ (.A1(_2666_),
    .A2(_2704_),
    .B(_2707_),
    .ZN(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7555_ (.A1(_2702_),
    .A2(_2703_),
    .B(_2708_),
    .ZN(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _7556_ (.A1(_2702_),
    .A2(_2703_),
    .A3(_2708_),
    .Z(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7557_ (.A1(_2709_),
    .A2(_2710_),
    .ZN(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7558_ (.A1(_2659_),
    .A2(_2711_),
    .ZN(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7559_ (.I(_2712_),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7560_ (.A1(_2701_),
    .A2(_2713_),
    .Z(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7561_ (.A1(_2694_),
    .A2(_2698_),
    .A3(_2714_),
    .Z(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7562_ (.A1(_2693_),
    .A2(_2715_),
    .Z(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7563_ (.A1(_2691_),
    .A2(_2716_),
    .Z(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7564_ (.I(_2718_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7565_ (.A1(_2646_),
    .A2(_2684_),
    .B(_2716_),
    .C(_2687_),
    .ZN(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7566_ (.A1(_2650_),
    .A2(_2681_),
    .B(_2693_),
    .ZN(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7567_ (.A1(_2682_),
    .A2(_2719_),
    .B1(_2720_),
    .B2(_2715_),
    .ZN(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7568_ (.A1(_2659_),
    .A2(_2711_),
    .B(_2709_),
    .ZN(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7569_ (.A1(_1688_),
    .A2(\C[1][16] ),
    .ZN(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7570_ (.A1(_1673_),
    .A2(_2707_),
    .A3(_2723_),
    .ZN(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7571_ (.A1(_2707_),
    .A2(_2723_),
    .B(_2724_),
    .ZN(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7572_ (.A1(_2722_),
    .A2(_2725_),
    .ZN(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7573_ (.A1(_2694_),
    .A2(_2714_),
    .Z(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7574_ (.A1(_2694_),
    .A2(_2714_),
    .Z(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7575_ (.A1(_2701_),
    .A2(_2713_),
    .B1(_2728_),
    .B2(_2698_),
    .C(_2729_),
    .ZN(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7576_ (.A1(_2721_),
    .A2(_2726_),
    .A3(_2730_),
    .Z(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7577_ (.I(_2731_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7578_ (.A1(_0048_),
    .A2(_0008_),
    .ZN(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _7579_ (.A1(_1597_),
    .A2(\C[0][0] ),
    .A3(_0757_),
    .A4(_0000_),
    .ZN(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7580_ (.A1(_1598_),
    .A2(\C[0][0] ),
    .A3(_1630_),
    .ZN(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7581_ (.A1(_0920_),
    .A2(_1772_),
    .B(_2734_),
    .ZN(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7582_ (.A1(_2733_),
    .A2(_2735_),
    .ZN(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7583_ (.A1(_2732_),
    .A2(_2736_),
    .Z(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7584_ (.I(_2738_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7585_ (.A1(_0209_),
    .A2(_0224_),
    .Z(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7586_ (.I(_2739_),
    .Z(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7587_ (.A1(_0950_),
    .A2(_0951_),
    .Z(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7588_ (.I(_2740_),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7589_ (.A1(_2732_),
    .A2(_2736_),
    .Z(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7590_ (.A1(_0033_),
    .A2(_1715_),
    .ZN(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7591_ (.A1(_0436_),
    .A2(_1826_),
    .ZN(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7592_ (.A1(_2742_),
    .A2(_2743_),
    .ZN(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7593_ (.A1(\C[0][1] ),
    .A2(_0184_),
    .ZN(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7594_ (.A1(_2744_),
    .A2(_2746_),
    .ZN(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7595_ (.A1(_2733_),
    .A2(_2747_),
    .ZN(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7596_ (.A1(_0375_),
    .A2(_1704_),
    .ZN(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7597_ (.A1(_0048_),
    .A2(_0009_),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7598_ (.A1(_2749_),
    .A2(_2750_),
    .Z(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7599_ (.A1(_2748_),
    .A2(_2751_),
    .ZN(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7600_ (.A1(_2741_),
    .A2(_2752_),
    .Z(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7601_ (.I(_2753_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7602_ (.A1(_0223_),
    .A2(_0225_),
    .Z(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7603_ (.I(_2754_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7604_ (.A1(_0944_),
    .A2(_0952_),
    .Z(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7605_ (.I(_2756_),
    .Z(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7606_ (.A1(_0375_),
    .A2(_1748_),
    .ZN(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7607_ (.A1(_0945_),
    .A2(_0010_),
    .B(_2757_),
    .ZN(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7608_ (.I(_0467_),
    .Z(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7609_ (.I(_2759_),
    .Z(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7610_ (.I(_2760_),
    .Z(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7611_ (.A1(_2761_),
    .A2(_0008_),
    .A3(_1759_),
    .A4(_2757_),
    .ZN(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7612_ (.A1(_0945_),
    .A2(_1704_),
    .A3(_0010_),
    .A4(_2757_),
    .ZN(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7613_ (.A1(_2762_),
    .A2(_2763_),
    .ZN(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7614_ (.A1(_2758_),
    .A2(_2765_),
    .ZN(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7615_ (.A1(_2733_),
    .A2(_2747_),
    .ZN(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7616_ (.A1(_2744_),
    .A2(_2746_),
    .ZN(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7617_ (.A1(_0897_),
    .A2(_1703_),
    .ZN(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7618_ (.A1(_2742_),
    .A2(_2743_),
    .Z(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7619_ (.I(_1713_),
    .Z(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7620_ (.A1(_0539_),
    .A2(_2771_),
    .ZN(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7621_ (.A1(_0922_),
    .A2(_0923_),
    .Z(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7622_ (.A1(_2773_),
    .A2(_1980_),
    .ZN(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7623_ (.A1(_0333_),
    .A2(net34),
    .ZN(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _7624_ (.A1(_2772_),
    .A2(_2774_),
    .A3(_2776_),
    .Z(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7625_ (.A1(\C[0][2] ),
    .A2(_0184_),
    .ZN(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7626_ (.A1(_2770_),
    .A2(_2777_),
    .A3(_2778_),
    .ZN(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7627_ (.A1(_2768_),
    .A2(_2769_),
    .A3(_2779_),
    .Z(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7628_ (.A1(_2767_),
    .A2(_2780_),
    .Z(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7629_ (.A1(_2766_),
    .A2(_2781_),
    .Z(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7630_ (.A1(_2748_),
    .A2(_2751_),
    .ZN(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7631_ (.A1(_2741_),
    .A2(_2752_),
    .ZN(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7632_ (.A1(_2783_),
    .A2(_2784_),
    .ZN(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7633_ (.A1(_2782_),
    .A2(_2785_),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7634_ (.I(_2787_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7635_ (.A1(_0230_),
    .A2(_0226_),
    .ZN(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7636_ (.A1(_0218_),
    .A2(_2788_),
    .ZN(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7637_ (.I(_2789_),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7638_ (.A1(_0940_),
    .A2(_0953_),
    .ZN(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7639_ (.A1(_0941_),
    .A2(_2790_),
    .ZN(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7640_ (.I(_2791_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7641_ (.A1(_2784_),
    .A2(_2782_),
    .ZN(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7642_ (.A1(_2783_),
    .A2(_2782_),
    .ZN(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7643_ (.A1(_2767_),
    .A2(_2780_),
    .Z(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7644_ (.A1(_2766_),
    .A2(_2781_),
    .B(_2795_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7645_ (.A1(_0375_),
    .A2(_1758_),
    .ZN(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7646_ (.A1(_2761_),
    .A2(_0011_),
    .B(_2797_),
    .ZN(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _7647_ (.A1(_2760_),
    .A2(_1762_),
    .A3(_1814_),
    .A4(_2797_),
    .ZN(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7648_ (.A1(_2761_),
    .A2(_1748_),
    .A3(_1812_),
    .A4(_2797_),
    .ZN(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7649_ (.A1(_2799_),
    .A2(_2800_),
    .ZN(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7650_ (.A1(_2798_),
    .A2(_2801_),
    .ZN(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7651_ (.A1(_2768_),
    .A2(_2779_),
    .ZN(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7652_ (.A1(_2768_),
    .A2(_2779_),
    .ZN(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7653_ (.A1(_0897_),
    .A2(_1704_),
    .A3(_2803_),
    .B(_2804_),
    .ZN(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7654_ (.A1(_2770_),
    .A2(_2777_),
    .ZN(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7655_ (.A1(_2807_),
    .A2(_2778_),
    .ZN(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7656_ (.A1(_2770_),
    .A2(_2777_),
    .ZN(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7657_ (.A1(_0752_),
    .A2(_1702_),
    .ZN(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7658_ (.A1(_0050_),
    .A2(_1762_),
    .A3(_2810_),
    .ZN(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7659_ (.A1(_0752_),
    .A2(_1703_),
    .B1(_1747_),
    .B2(_0896_),
    .ZN(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7660_ (.A1(_2811_),
    .A2(_2812_),
    .ZN(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7661_ (.A1(_2809_),
    .A2(_2813_),
    .ZN(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7662_ (.A1(_0348_),
    .A2(_0352_),
    .Z(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7663_ (.A1(_2815_),
    .A2(_1771_),
    .B1(_1972_),
    .B2(_2773_),
    .ZN(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7664_ (.A1(_2815_),
    .A2(_2773_),
    .A3(_1771_),
    .A4(_1972_),
    .ZN(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7665_ (.A1(_2817_),
    .A2(_2776_),
    .B(_2818_),
    .ZN(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7666_ (.A1(_0823_),
    .A2(_1783_),
    .ZN(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7667_ (.A1(_0924_),
    .A2(_1975_),
    .ZN(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7668_ (.A1(_0435_),
    .A2(_0003_),
    .ZN(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7669_ (.A1(_2820_),
    .A2(_2821_),
    .A3(_2822_),
    .Z(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7670_ (.I(_0403_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7671_ (.A1(_1479_),
    .A2(\C[0][3] ),
    .Z(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7672_ (.A1(_0035_),
    .A2(_1716_),
    .A3(_2824_),
    .Z(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7673_ (.A1(_0035_),
    .A2(_1716_),
    .B1(_2824_),
    .B2(_1534_),
    .ZN(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7674_ (.A1(_2825_),
    .A2(_2827_),
    .ZN(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7675_ (.A1(_2819_),
    .A2(_2823_),
    .A3(_2828_),
    .ZN(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7676_ (.A1(_2808_),
    .A2(_2814_),
    .A3(_2829_),
    .ZN(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7677_ (.A1(_2802_),
    .A2(_2806_),
    .A3(_2830_),
    .ZN(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7678_ (.A1(_2762_),
    .A2(_2796_),
    .A3(_2831_),
    .ZN(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7679_ (.A1(_2793_),
    .A2(_2832_),
    .Z(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7680_ (.A1(_2792_),
    .A2(_2833_),
    .Z(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7681_ (.I(_2834_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7682_ (.A1(_0228_),
    .A2(_0254_),
    .Z(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7683_ (.I(_2835_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7684_ (.A1(_0954_),
    .A2(_0955_),
    .Z(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7685_ (.I(_2837_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7686_ (.A1(_2783_),
    .A2(_2782_),
    .A3(_2832_),
    .ZN(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _7687_ (.A1(_2792_),
    .A2(_2833_),
    .B(_2838_),
    .ZN(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7688_ (.A1(_2796_),
    .A2(_2831_),
    .Z(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7689_ (.A1(_2796_),
    .A2(_2831_),
    .Z(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7690_ (.A1(_2762_),
    .A2(_2840_),
    .B(_2841_),
    .ZN(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7691_ (.A1(_2806_),
    .A2(_2830_),
    .ZN(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7692_ (.A1(_2806_),
    .A2(_2830_),
    .ZN(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7693_ (.A1(_2798_),
    .A2(_2801_),
    .A3(_2843_),
    .B(_2844_),
    .ZN(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7694_ (.A1(_0945_),
    .A2(_0011_),
    .A3(_2797_),
    .ZN(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7695_ (.A1(_2770_),
    .A2(_2777_),
    .A3(_2813_),
    .ZN(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7696_ (.A1(_0903_),
    .A2(_1811_),
    .ZN(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7697_ (.A1(_2849_),
    .A2(_2811_),
    .Z(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7698_ (.A1(_2759_),
    .A2(_1865_),
    .ZN(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7699_ (.A1(_2850_),
    .A2(_2851_),
    .ZN(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7700_ (.A1(_2848_),
    .A2(_2852_),
    .Z(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7701_ (.A1(_2847_),
    .A2(_2853_),
    .Z(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7702_ (.A1(_2807_),
    .A2(_2778_),
    .B(_2829_),
    .ZN(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7703_ (.A1(_2807_),
    .A2(_2778_),
    .A3(_2829_),
    .ZN(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7704_ (.A1(_2814_),
    .A2(_2855_),
    .B(_2857_),
    .ZN(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7705_ (.A1(_2819_),
    .A2(_2823_),
    .Z(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7706_ (.A1(_2819_),
    .A2(_2823_),
    .ZN(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _7707_ (.A1(_2859_),
    .A2(_2860_),
    .A3(_2825_),
    .A4(_2827_),
    .ZN(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7708_ (.A1(_0751_),
    .A2(_1746_),
    .ZN(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7709_ (.A1(_0761_),
    .A2(_1701_),
    .ZN(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7710_ (.A1(_0335_),
    .A2(_0896_),
    .A3(_2237_),
    .ZN(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7711_ (.A1(_2862_),
    .A2(_2863_),
    .A3(_2864_),
    .Z(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7712_ (.A1(_2860_),
    .A2(_2865_),
    .Z(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7713_ (.A1(_0899_),
    .A2(_0001_),
    .B1(_0002_),
    .B2(_0925_),
    .ZN(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7714_ (.A1(_0034_),
    .A2(_0925_),
    .A3(_1736_),
    .A4(_0002_),
    .ZN(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7715_ (.A1(_2868_),
    .A2(_2822_),
    .B(_2869_),
    .ZN(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7716_ (.A1(_3037_),
    .A2(_1731_),
    .B(\A[0][2] ),
    .ZN(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _7717_ (.A1(_2826_),
    .A2(_1848_),
    .ZN(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7718_ (.A1(_0348_),
    .A2(_0352_),
    .B1(_2871_),
    .B2(_2872_),
    .C(_2236_),
    .ZN(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7719_ (.A1(_0922_),
    .A2(_0923_),
    .B1(_1847_),
    .B2(_1850_),
    .C(_4066_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7720_ (.A1(_2873_),
    .A2(_2874_),
    .Z(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7721_ (.A1(_0334_),
    .A2(_1999_),
    .ZN(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7722_ (.A1(_2875_),
    .A2(_2876_),
    .Z(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7723_ (.A1(_2870_),
    .A2(_2877_),
    .Z(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7724_ (.A1(_0035_),
    .A2(_1716_),
    .A3(_2824_),
    .ZN(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7725_ (.A1(_0488_),
    .A2(_2771_),
    .ZN(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7726_ (.A1(_0775_),
    .A2(_1783_),
    .ZN(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7727_ (.A1(\C[0][4] ),
    .A2(_4239_),
    .ZN(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7728_ (.A1(_2881_),
    .A2(_2882_),
    .A3(_2883_),
    .Z(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7729_ (.A1(_2880_),
    .A2(_2884_),
    .Z(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7730_ (.A1(_2879_),
    .A2(_2885_),
    .Z(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7731_ (.A1(_2861_),
    .A2(_2866_),
    .A3(_2886_),
    .ZN(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7732_ (.A1(_2858_),
    .A2(_2887_),
    .ZN(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7733_ (.A1(_2854_),
    .A2(_2888_),
    .Z(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7734_ (.A1(_2799_),
    .A2(_2846_),
    .A3(_2890_),
    .ZN(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7735_ (.A1(_2842_),
    .A2(_2891_),
    .Z(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7736_ (.A1(_2839_),
    .A2(_2892_),
    .Z(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7737_ (.I(_2893_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7738_ (.A1(_0259_),
    .A2(_0275_),
    .A3(_0256_),
    .ZN(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7739_ (.I(_2894_),
    .Z(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7740_ (.A1(_0956_),
    .A2(_0957_),
    .Z(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7741_ (.I(_2895_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7742_ (.A1(_2842_),
    .A2(_2891_),
    .Z(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7743_ (.A1(_2839_),
    .A2(_2892_),
    .B(_2896_),
    .ZN(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7744_ (.A1(_2846_),
    .A2(_2890_),
    .ZN(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7745_ (.A1(_2846_),
    .A2(_2890_),
    .ZN(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7746_ (.A1(_2799_),
    .A2(_2899_),
    .B(_2900_),
    .ZN(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7747_ (.A1(_2848_),
    .A2(_2852_),
    .ZN(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7748_ (.A1(_2848_),
    .A2(_2852_),
    .ZN(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7749_ (.A1(_2847_),
    .A2(_2902_),
    .B(_2903_),
    .ZN(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7750_ (.A1(_2858_),
    .A2(_2887_),
    .Z(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7751_ (.A1(_2854_),
    .A2(_2888_),
    .B(_2905_),
    .ZN(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7752_ (.A1(_2761_),
    .A2(_0012_),
    .A3(_2850_),
    .ZN(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7753_ (.A1(_2849_),
    .A2(_2811_),
    .B(_2907_),
    .ZN(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7754_ (.A1(_2860_),
    .A2(_2865_),
    .Z(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7755_ (.I(_1744_),
    .Z(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7756_ (.A1(_4158_),
    .A2(_0761_),
    .A3(_2911_),
    .ZN(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7757_ (.A1(_0335_),
    .A2(_0752_),
    .A3(_2911_),
    .B1(_1702_),
    .B2(_0761_),
    .ZN(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7758_ (.A1(_2810_),
    .A2(_2912_),
    .B1(_2913_),
    .B2(_2864_),
    .ZN(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7759_ (.A1(_0838_),
    .A2(_2120_),
    .ZN(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7760_ (.A1(_2914_),
    .A2(_2915_),
    .Z(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7761_ (.A1(_2759_),
    .A2(_1931_),
    .Z(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7762_ (.A1(_2916_),
    .A2(_2917_),
    .Z(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7763_ (.A1(_2910_),
    .A2(_2918_),
    .Z(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7764_ (.A1(_2909_),
    .A2(_2920_),
    .Z(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7765_ (.A1(_2861_),
    .A2(_2886_),
    .Z(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7766_ (.A1(_2861_),
    .A2(_2886_),
    .Z(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7767_ (.A1(_2866_),
    .A2(_2922_),
    .B(_2923_),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7768_ (.A1(_2870_),
    .A2(_2877_),
    .ZN(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7769_ (.A1(_0308_),
    .A2(_1701_),
    .ZN(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7770_ (.A1(_0896_),
    .A2(_1814_),
    .ZN(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7771_ (.A1(_4158_),
    .A2(_0751_),
    .A3(_2237_),
    .ZN(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7772_ (.A1(_2912_),
    .A2(_2928_),
    .Z(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7773_ (.A1(_2927_),
    .A2(_2929_),
    .Z(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7774_ (.A1(_2926_),
    .A2(_2931_),
    .ZN(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7775_ (.A1(_2925_),
    .A2(_2932_),
    .ZN(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7776_ (.A1(_2880_),
    .A2(_2884_),
    .ZN(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7777_ (.A1(_2879_),
    .A2(_2885_),
    .B(_2934_),
    .ZN(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7778_ (.A1(_2873_),
    .A2(_2874_),
    .Z(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7779_ (.A1(_2875_),
    .A2(_2876_),
    .B(_2936_),
    .ZN(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _7780_ (.A1(_0391_),
    .A2(_0400_),
    .A3(_1713_),
    .A4(_1735_),
    .ZN(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7781_ (.A1(_0348_),
    .A2(_0352_),
    .B1(_1847_),
    .B2(_1850_),
    .C(_3593_),
    .ZN(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7782_ (.A1(_0922_),
    .A2(_0923_),
    .B1(_1897_),
    .B2(_1898_),
    .C(_3991_),
    .ZN(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7783_ (.A1(_2939_),
    .A2(_2940_),
    .Z(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7784_ (.A1(_0435_),
    .A2(_2257_),
    .Z(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7785_ (.A1(_2938_),
    .A2(_2942_),
    .A3(_2943_),
    .Z(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7786_ (.A1(_2937_),
    .A2(_2944_),
    .ZN(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7787_ (.A1(_0379_),
    .A2(_0381_),
    .Z(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7788_ (.A1(_0387_),
    .A2(_0388_),
    .Z(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7789_ (.A1(_2946_),
    .A2(_1771_),
    .B1(_1972_),
    .B2(_2947_),
    .ZN(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7790_ (.A1(\C[0][4] ),
    .A2(_3929_),
    .A3(_2938_),
    .A4(_2948_),
    .ZN(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7791_ (.A1(_0571_),
    .A2(_1714_),
    .ZN(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7792_ (.A1(_0383_),
    .A2(net38),
    .ZN(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7793_ (.A1(_0389_),
    .A2(_1894_),
    .ZN(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7794_ (.A1(_2950_),
    .A2(_2951_),
    .A3(_2953_),
    .Z(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7795_ (.A1(\C[0][5] ),
    .A2(_4239_),
    .ZN(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7796_ (.I(_2955_),
    .Z(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _7797_ (.A1(_2949_),
    .A2(_2954_),
    .A3(_2956_),
    .Z(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7798_ (.A1(_2945_),
    .A2(_2957_),
    .Z(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7799_ (.A1(_2935_),
    .A2(_2958_),
    .Z(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7800_ (.A1(_2933_),
    .A2(_2959_),
    .ZN(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7801_ (.A1(_2921_),
    .A2(_2924_),
    .A3(_2960_),
    .Z(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7802_ (.A1(_2906_),
    .A2(_2961_),
    .Z(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7803_ (.A1(_2904_),
    .A2(_2962_),
    .Z(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7804_ (.A1(_2898_),
    .A2(_2901_),
    .A3(_2964_),
    .ZN(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7805_ (.I(_2965_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7806_ (.A1(_0278_),
    .A2(_0291_),
    .Z(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7807_ (.I(_2966_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7808_ (.A1(_0934_),
    .A2(_0958_),
    .ZN(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7809_ (.A1(_2967_),
    .A2(_0959_),
    .ZN(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7810_ (.I(_2968_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7811_ (.A1(_2906_),
    .A2(_2961_),
    .Z(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7812_ (.A1(_2904_),
    .A2(_2962_),
    .B(_2969_),
    .ZN(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7813_ (.A1(_2910_),
    .A2(_2918_),
    .ZN(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7814_ (.A1(_2909_),
    .A2(_2920_),
    .ZN(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7815_ (.A1(_2972_),
    .A2(_2973_),
    .ZN(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7816_ (.A1(_2924_),
    .A2(_2960_),
    .ZN(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7817_ (.A1(_2924_),
    .A2(_2960_),
    .ZN(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7818_ (.A1(_2921_),
    .A2(_2975_),
    .B(_2976_),
    .ZN(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7819_ (.A1(_2914_),
    .A2(_2915_),
    .ZN(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7820_ (.A1(_2916_),
    .A2(_2917_),
    .B(_2978_),
    .ZN(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7821_ (.A1(_2925_),
    .A2(_2932_),
    .Z(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7822_ (.A1(_1753_),
    .A2(_0317_),
    .A3(_1755_),
    .ZN(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7823_ (.A1(_2862_),
    .A2(_2981_),
    .B1(_2929_),
    .B2(_2927_),
    .ZN(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7824_ (.A1(_0838_),
    .A2(_1952_),
    .ZN(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7825_ (.A1(_2983_),
    .A2(_2984_),
    .ZN(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7826_ (.A1(_2759_),
    .A2(_2014_),
    .ZN(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7827_ (.A1(_2985_),
    .A2(_2986_),
    .ZN(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7828_ (.A1(_2980_),
    .A2(_2987_),
    .ZN(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7829_ (.A1(_2979_),
    .A2(_2988_),
    .ZN(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7830_ (.A1(_2879_),
    .A2(_2885_),
    .Z(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7831_ (.A1(_2934_),
    .A2(_2990_),
    .B(_2958_),
    .ZN(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7832_ (.A1(_2933_),
    .A2(_2959_),
    .B(_2991_),
    .ZN(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7833_ (.A1(_2926_),
    .A2(_2931_),
    .ZN(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7834_ (.A1(_2942_),
    .A2(_2943_),
    .Z(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7835_ (.A1(_2942_),
    .A2(_2943_),
    .ZN(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7836_ (.A1(_2938_),
    .A2(_2995_),
    .A3(_2996_),
    .B1(_2944_),
    .B2(_2937_),
    .ZN(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7837_ (.A1(_0326_),
    .A2(_1823_),
    .ZN(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7838_ (.A1(_2236_),
    .A2(_0307_),
    .A3(_2911_),
    .ZN(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7839_ (.A1(_2998_),
    .A2(_2999_),
    .ZN(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7840_ (.A1(_0344_),
    .A2(_1863_),
    .ZN(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7841_ (.I(_1807_),
    .Z(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7842_ (.A1(_3793_),
    .A2(_0751_),
    .A3(_3002_),
    .ZN(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7843_ (.A1(_2981_),
    .A2(_3001_),
    .A3(_3003_),
    .ZN(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7844_ (.A1(_3000_),
    .A2(_3005_),
    .ZN(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7845_ (.A1(_2997_),
    .A2(_3006_),
    .ZN(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7846_ (.A1(_2994_),
    .A2(_3007_),
    .ZN(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7847_ (.I(_2954_),
    .Z(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7848_ (.A1(_3009_),
    .A2(_2956_),
    .ZN(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7849_ (.A1(_3009_),
    .A2(_2956_),
    .Z(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _7850_ (.A1(_2949_),
    .A2(_3010_),
    .A3(_3011_),
    .B1(_2957_),
    .B2(_2945_),
    .ZN(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7851_ (.A1(_0479_),
    .A2(_0480_),
    .B1(_1732_),
    .B2(_1734_),
    .C(_2867_),
    .ZN(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7852_ (.A1(_0379_),
    .A2(_0381_),
    .B1(_2871_),
    .B2(_2872_),
    .C(_3100_),
    .ZN(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _7853_ (.A1(_0387_),
    .A2(_0388_),
    .B1(_1847_),
    .B2(_1850_),
    .C(_1753_),
    .ZN(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7854_ (.A1(_3013_),
    .A2(_3014_),
    .A3(_3016_),
    .Z(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _7855_ (.A1(_0514_),
    .A2(\C[0][6] ),
    .A3(_0569_),
    .A4(net43),
    .ZN(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7856_ (.A1(_0504_),
    .A2(_0505_),
    .Z(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7857_ (.A1(_0473_),
    .A2(\C[0][6] ),
    .ZN(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7858_ (.A1(_3019_),
    .A2(_1770_),
    .B1(_3020_),
    .B2(_1181_),
    .ZN(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7859_ (.A1(_3017_),
    .A2(_3018_),
    .A3(_3021_),
    .Z(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7860_ (.I(_3022_),
    .Z(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7861_ (.A1(_3018_),
    .A2(_3021_),
    .B(_3017_),
    .ZN(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7862_ (.A1(_3023_),
    .A2(_3024_),
    .ZN(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7863_ (.A1(_2939_),
    .A2(_2940_),
    .Z(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7864_ (.A1(_2942_),
    .A2(_2943_),
    .B(_3027_),
    .ZN(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7865_ (.A1(_0720_),
    .A2(_2771_),
    .B1(_1781_),
    .B2(_0383_),
    .ZN(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7866_ (.A1(_0401_),
    .A2(_1252_),
    .A3(_1714_),
    .A4(_1736_),
    .ZN(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7867_ (.A1(_3029_),
    .A2(_2953_),
    .B(_3030_),
    .ZN(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7868_ (.A1(_0822_),
    .A2(_2055_),
    .ZN(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7869_ (.A1(_0924_),
    .A2(_2257_),
    .ZN(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7870_ (.A1(_0435_),
    .A2(_2562_),
    .ZN(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7871_ (.A1(_3032_),
    .A2(_3033_),
    .A3(_3034_),
    .ZN(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7872_ (.A1(_3028_),
    .A2(_3031_),
    .A3(_3035_),
    .ZN(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7873_ (.A1(_3010_),
    .A2(_3025_),
    .A3(_3036_),
    .Z(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7874_ (.A1(_3008_),
    .A2(_3012_),
    .A3(_3038_),
    .ZN(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7875_ (.A1(_2992_),
    .A2(_3039_),
    .ZN(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7876_ (.A1(_2989_),
    .A2(_3040_),
    .Z(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _7877_ (.A1(_2974_),
    .A2(_2977_),
    .A3(_3041_),
    .Z(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7878_ (.A1(_2970_),
    .A2(_3042_),
    .ZN(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7879_ (.A1(_2901_),
    .A2(_2964_),
    .ZN(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7880_ (.A1(_2839_),
    .A2(_2892_),
    .B1(_2901_),
    .B2(_2964_),
    .C(_2896_),
    .ZN(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7881_ (.A1(_3044_),
    .A2(_3045_),
    .ZN(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7882_ (.A1(_3043_),
    .A2(_3046_),
    .ZN(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7883_ (.I(_3047_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7884_ (.A1(_0293_),
    .A2(_0298_),
    .Z(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7885_ (.I(_3049_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7886_ (.A1(_0918_),
    .A2(_0960_),
    .ZN(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7887_ (.A1(_3050_),
    .A2(_0961_),
    .ZN(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7888_ (.I(_3051_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _7889_ (.A1(_3044_),
    .A2(_3043_),
    .A3(_3045_),
    .B1(_2970_),
    .B2(_3042_),
    .ZN(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7890_ (.I(_2977_),
    .ZN(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7891_ (.A1(_3053_),
    .A2(_3041_),
    .ZN(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7892_ (.A1(_2977_),
    .A2(_3041_),
    .ZN(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7893_ (.A1(_2974_),
    .A2(_3055_),
    .ZN(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7894_ (.A1(_2980_),
    .A2(_2987_),
    .ZN(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7895_ (.A1(_2979_),
    .A2(_2988_),
    .ZN(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7896_ (.A1(_3058_),
    .A2(_3059_),
    .ZN(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7897_ (.A1(_2992_),
    .A2(_3039_),
    .ZN(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7898_ (.A1(_2989_),
    .A2(_3040_),
    .B(_3061_),
    .ZN(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7899_ (.A1(_2983_),
    .A2(_2984_),
    .Z(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7900_ (.A1(_2985_),
    .A2(_2986_),
    .B(_3063_),
    .ZN(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7901_ (.A1(_2997_),
    .A2(_3006_),
    .ZN(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7902_ (.A1(_2994_),
    .A2(_3007_),
    .B(_3065_),
    .ZN(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7903_ (.A1(_2981_),
    .A2(_3003_),
    .ZN(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7904_ (.A1(_3792_),
    .A2(_0317_),
    .A3(_3002_),
    .ZN(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7905_ (.A1(_2928_),
    .A2(_3069_),
    .ZN(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7906_ (.A1(_3001_),
    .A2(_3068_),
    .B(_3070_),
    .ZN(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7907_ (.A1(_0903_),
    .A2(_2579_),
    .ZN(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7908_ (.A1(_3071_),
    .A2(_3072_),
    .ZN(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7909_ (.A1(_2760_),
    .A2(_2203_),
    .ZN(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7910_ (.A1(_3073_),
    .A2(_3074_),
    .ZN(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7911_ (.A1(_3066_),
    .A2(_3075_),
    .Z(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7912_ (.A1(_3064_),
    .A2(_3076_),
    .ZN(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7913_ (.A1(_3012_),
    .A2(_3038_),
    .ZN(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7914_ (.A1(_3012_),
    .A2(_3038_),
    .ZN(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7915_ (.A1(_3008_),
    .A2(_3079_),
    .B(_3080_),
    .ZN(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7916_ (.I(_3005_),
    .ZN(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7917_ (.A1(_3000_),
    .A2(_3082_),
    .ZN(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7918_ (.A1(_3027_),
    .A2(_2995_),
    .Z(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7919_ (.A1(_3031_),
    .A2(_3035_),
    .Z(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7920_ (.A1(_3031_),
    .A2(_3035_),
    .Z(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7921_ (.A1(_3084_),
    .A2(_3085_),
    .B(_3086_),
    .ZN(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7922_ (.A1(_3960_),
    .A2(_0325_),
    .A3(_2050_),
    .ZN(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7923_ (.A1(_2926_),
    .A2(_3088_),
    .Z(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7924_ (.A1(_0363_),
    .A2(_1929_),
    .ZN(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7925_ (.A1(_0314_),
    .A2(_1862_),
    .ZN(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7926_ (.A1(_3069_),
    .A2(_3092_),
    .ZN(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7927_ (.A1(_3091_),
    .A2(_3093_),
    .ZN(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7928_ (.A1(_3992_),
    .A2(_0307_),
    .A3(_2237_),
    .ZN(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7929_ (.A1(_0577_),
    .A2(_1823_),
    .ZN(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7930_ (.A1(_3088_),
    .A2(_3095_),
    .A3(_3096_),
    .Z(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _7931_ (.A1(_3090_),
    .A2(_3094_),
    .A3(_3097_),
    .ZN(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7932_ (.A1(_3083_),
    .A2(_3087_),
    .A3(_3098_),
    .ZN(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7933_ (.A1(_3009_),
    .A2(_2956_),
    .B1(_3023_),
    .B2(_3024_),
    .ZN(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7934_ (.A1(_3009_),
    .A2(_2955_),
    .A3(_3023_),
    .A4(_3024_),
    .ZN(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7935_ (.A1(_3101_),
    .A2(_3036_),
    .B(_3102_),
    .ZN(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7936_ (.A1(_2871_),
    .A2(_2872_),
    .ZN(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7937_ (.A1(_0382_),
    .A2(_0509_),
    .A3(_3104_),
    .A4(_2275_),
    .Z(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7938_ (.A1(_0481_),
    .A2(_1841_),
    .B1(_1903_),
    .B2(_0382_),
    .ZN(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7939_ (.A1(_3105_),
    .A2(_3106_),
    .Z(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7940_ (.A1(_0392_),
    .A2(_2250_),
    .ZN(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7941_ (.A1(_3107_),
    .A2(_3108_),
    .Z(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7942_ (.I(\C[0][7] ),
    .ZN(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7943_ (.A1(_3423_),
    .A2(_3110_),
    .ZN(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7944_ (.A1(_0651_),
    .A2(_1714_),
    .A3(_3112_),
    .ZN(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7945_ (.A1(_3434_),
    .A2(_3110_),
    .A3(_1181_),
    .B1(_0566_),
    .B2(_1770_),
    .ZN(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7946_ (.A1(_3113_),
    .A2(_3114_),
    .ZN(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7947_ (.A1(_3019_),
    .A2(_1980_),
    .ZN(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7948_ (.A1(_3018_),
    .A2(_3115_),
    .A3(_3116_),
    .Z(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7949_ (.A1(_3023_),
    .A2(_3109_),
    .A3(_3117_),
    .Z(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7950_ (.A1(_3032_),
    .A2(_3033_),
    .Z(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7951_ (.A1(_3032_),
    .A2(_3033_),
    .Z(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7952_ (.A1(_3119_),
    .A2(_3034_),
    .B(_3120_),
    .ZN(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7953_ (.A1(_3013_),
    .A2(_3014_),
    .ZN(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7954_ (.A1(_0389_),
    .A2(_1962_),
    .ZN(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7955_ (.A1(_3013_),
    .A2(_3014_),
    .ZN(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7956_ (.A1(_3123_),
    .A2(_3124_),
    .B(_3125_),
    .ZN(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7957_ (.A1(_0822_),
    .A2(_2185_),
    .ZN(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7958_ (.A1(_0360_),
    .A2(_2077_),
    .ZN(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7959_ (.A1(_0434_),
    .A2(_2281_),
    .Z(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7960_ (.A1(_3127_),
    .A2(_3128_),
    .A3(_3129_),
    .Z(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7961_ (.A1(_3126_),
    .A2(_3130_),
    .Z(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7962_ (.A1(_3121_),
    .A2(_3131_),
    .Z(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7963_ (.A1(_3103_),
    .A2(_3118_),
    .A3(_3132_),
    .Z(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7964_ (.A1(_3099_),
    .A2(_3134_),
    .Z(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7965_ (.A1(_3081_),
    .A2(_3135_),
    .ZN(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7966_ (.A1(_3077_),
    .A2(_3136_),
    .Z(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7967_ (.A1(_3062_),
    .A2(_3137_),
    .ZN(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7968_ (.A1(_3060_),
    .A2(_3138_),
    .ZN(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7969_ (.A1(_3054_),
    .A2(_3057_),
    .A3(_3139_),
    .ZN(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7970_ (.A1(_3054_),
    .A2(_3057_),
    .B(_3139_),
    .ZN(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7971_ (.I(_3141_),
    .ZN(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7972_ (.A1(_3140_),
    .A2(_3142_),
    .ZN(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7973_ (.A1(_3052_),
    .A2(_3143_),
    .ZN(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7974_ (.I(_3145_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7975_ (.A1(_0293_),
    .A2(_0298_),
    .B(_0299_),
    .ZN(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7976_ (.A1(_0176_),
    .A2(_0177_),
    .A3(_3146_),
    .Z(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7977_ (.I(_3147_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7978_ (.A1(_0893_),
    .A2(_0962_),
    .ZN(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7979_ (.A1(_3148_),
    .A2(_0963_),
    .ZN(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7980_ (.I(_3149_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7981_ (.A1(_3066_),
    .A2(_3075_),
    .ZN(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7982_ (.A1(_3064_),
    .A2(_3076_),
    .ZN(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7983_ (.A1(_3150_),
    .A2(_3151_),
    .ZN(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7984_ (.A1(_3081_),
    .A2(_3135_),
    .ZN(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7985_ (.A1(_3077_),
    .A2(_3136_),
    .B(_3154_),
    .ZN(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7986_ (.A1(_0049_),
    .A2(_0014_),
    .A3(_3071_),
    .ZN(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7987_ (.A1(_2760_),
    .A2(_2103_),
    .A3(_3073_),
    .ZN(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7988_ (.A1(_3156_),
    .A2(_3157_),
    .ZN(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7989_ (.A1(_3087_),
    .A2(_3098_),
    .ZN(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _7990_ (.A1(_3000_),
    .A2(_3082_),
    .A3(_3159_),
    .B1(_3098_),
    .B2(_3087_),
    .ZN(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7991_ (.A1(_0052_),
    .A2(_1865_),
    .A3(_3003_),
    .ZN(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7992_ (.A1(_0050_),
    .A2(_0013_),
    .A3(_3093_),
    .ZN(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7993_ (.A1(_3161_),
    .A2(_3162_),
    .ZN(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7994_ (.A1(_0049_),
    .A2(_2203_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7995_ (.A1(_3164_),
    .A2(_3165_),
    .ZN(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7996_ (.A1(_3158_),
    .A2(_3160_),
    .A3(_3166_),
    .ZN(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7997_ (.I(_3022_),
    .ZN(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7998_ (.A1(_3168_),
    .A2(_3109_),
    .A3(_3117_),
    .Z(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7999_ (.A1(_3121_),
    .A2(_3131_),
    .ZN(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8000_ (.A1(_3169_),
    .A2(_3170_),
    .ZN(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8001_ (.A1(_3118_),
    .A2(_3132_),
    .ZN(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _8002_ (.A1(_3103_),
    .A2(_3171_),
    .A3(_3172_),
    .B1(_3134_),
    .B2(_3099_),
    .ZN(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8003_ (.A1(_3090_),
    .A2(_3097_),
    .Z(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8004_ (.A1(_3090_),
    .A2(_3097_),
    .Z(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8005_ (.A1(_3094_),
    .A2(_3175_),
    .B(_3176_),
    .ZN(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8006_ (.A1(_3126_),
    .A2(_3130_),
    .Z(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _8007_ (.A1(_3121_),
    .A2(_3131_),
    .B(_3178_),
    .ZN(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8008_ (.A1(_0413_),
    .A2(_2012_),
    .ZN(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8009_ (.A1(_0319_),
    .A2(_2045_),
    .ZN(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8010_ (.A1(_0529_),
    .A2(_1928_),
    .ZN(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8011_ (.A1(_3181_),
    .A2(_3182_),
    .ZN(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8012_ (.A1(_3180_),
    .A2(_3183_),
    .ZN(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8013_ (.A1(_3947_),
    .A2(_0576_),
    .A3(_2050_),
    .ZN(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _8014_ (.A1(_1184_),
    .A2(_0326_),
    .A3(_2911_),
    .B1(_1701_),
    .B2(_0577_),
    .ZN(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8015_ (.A1(_2998_),
    .A2(_3186_),
    .B1(_3187_),
    .B2(_3095_),
    .ZN(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8016_ (.A1(_3947_),
    .A2(_0325_),
    .A3(_1755_),
    .ZN(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8017_ (.A1(_2236_),
    .A2(_0308_),
    .A3(_3002_),
    .ZN(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8018_ (.A1(_3186_),
    .A2(_3189_),
    .A3(_3190_),
    .Z(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8019_ (.A1(_3188_),
    .A2(_3191_),
    .Z(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8020_ (.A1(_3184_),
    .A2(_3192_),
    .Z(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _8021_ (.A1(_3177_),
    .A2(_3179_),
    .A3(_3193_),
    .ZN(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8022_ (.A1(_3109_),
    .A2(_3117_),
    .Z(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8023_ (.A1(_3109_),
    .A2(_3117_),
    .ZN(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _8024_ (.A1(_3168_),
    .A2(_3195_),
    .A3(_3197_),
    .B1(_3169_),
    .B2(_3170_),
    .ZN(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8025_ (.A1(_3127_),
    .A2(_3128_),
    .ZN(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8026_ (.A1(_3127_),
    .A2(_3128_),
    .ZN(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8027_ (.A1(_3199_),
    .A2(_3129_),
    .B(_3200_),
    .ZN(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8028_ (.A1(_0384_),
    .A2(_1252_),
    .A3(_3104_),
    .A4(_1907_),
    .ZN(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8029_ (.A1(_3106_),
    .A2(_3108_),
    .B(_3202_),
    .ZN(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8030_ (.A1(_0822_),
    .A2(_2350_),
    .ZN(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8031_ (.A1(_0924_),
    .A2(_2404_),
    .ZN(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8032_ (.A1(_3204_),
    .A2(_3205_),
    .Z(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8033_ (.A1(_3201_),
    .A2(_3203_),
    .A3(_3206_),
    .Z(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8034_ (.A1(_3107_),
    .A2(_3108_),
    .ZN(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8035_ (.A1(_3113_),
    .A2(_3114_),
    .A3(_3116_),
    .ZN(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _8036_ (.A1(_0716_),
    .A2(_1715_),
    .A3(_3112_),
    .Z(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8037_ (.A1(_0716_),
    .A2(_2771_),
    .B1(_3112_),
    .B2(_3976_),
    .ZN(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8038_ (.A1(_0718_),
    .A2(_1736_),
    .ZN(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8039_ (.A1(_3211_),
    .A2(_3212_),
    .B(_3213_),
    .ZN(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8040_ (.I(_3018_),
    .ZN(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8041_ (.A1(_3210_),
    .A2(_3214_),
    .B(_3215_),
    .ZN(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8042_ (.A1(_3215_),
    .A2(_3210_),
    .A3(_3214_),
    .ZN(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8043_ (.A1(_3209_),
    .A2(_3216_),
    .B(_3217_),
    .ZN(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8044_ (.A1(_0403_),
    .A2(_1987_),
    .ZN(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8045_ (.A1(_1252_),
    .A2(_1851_),
    .ZN(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8046_ (.A1(_0487_),
    .A2(_2250_),
    .ZN(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8047_ (.A1(_3221_),
    .A2(_3222_),
    .ZN(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8048_ (.A1(_3220_),
    .A2(_3223_),
    .Z(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8049_ (.A1(_3212_),
    .A2(_3213_),
    .B(_3113_),
    .ZN(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8050_ (.A1(_0456_),
    .A2(\C[0][8] ),
    .ZN(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8051_ (.A1(_3926_),
    .A2(_3226_),
    .ZN(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _8052_ (.A1(_0564_),
    .A2(_0565_),
    .B1(_1732_),
    .B2(_1734_),
    .C(_3960_),
    .ZN(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8053_ (.I0(_3227_),
    .I1(_3226_),
    .S(_3228_),
    .Z(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8054_ (.A1(_0633_),
    .A2(_3104_),
    .ZN(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8055_ (.A1(_3230_),
    .A2(_3231_),
    .ZN(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8056_ (.A1(_3225_),
    .A2(_3232_),
    .Z(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8057_ (.A1(_3224_),
    .A2(_3233_),
    .Z(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _8058_ (.A1(_3208_),
    .A2(_3219_),
    .A3(_3234_),
    .ZN(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8059_ (.A1(_3194_),
    .A2(_3198_),
    .A3(_3235_),
    .Z(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8060_ (.A1(_3173_),
    .A2(_3236_),
    .Z(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8061_ (.A1(_3167_),
    .A2(_3237_),
    .ZN(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8062_ (.A1(_3155_),
    .A2(_3238_),
    .ZN(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8063_ (.A1(_3153_),
    .A2(_3239_),
    .ZN(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8064_ (.A1(_3062_),
    .A2(_3137_),
    .ZN(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8065_ (.A1(_3060_),
    .A2(_3138_),
    .B(_3242_),
    .ZN(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8066_ (.A1(_3241_),
    .A2(_3243_),
    .ZN(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8067_ (.A1(_3052_),
    .A2(_3140_),
    .ZN(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8068_ (.A1(_3142_),
    .A2(_3245_),
    .ZN(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8069_ (.A1(_3244_),
    .A2(_3246_),
    .Z(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8070_ (.I(_3247_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8071_ (.A1(_0965_),
    .A2(_0967_),
    .Z(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8072_ (.I(_3248_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8073_ (.I(_3238_),
    .ZN(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8074_ (.A1(_3155_),
    .A2(_3250_),
    .ZN(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8075_ (.A1(_3153_),
    .A2(_3239_),
    .ZN(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8076_ (.A1(_3251_),
    .A2(_3252_),
    .ZN(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8077_ (.A1(_3160_),
    .A2(_3166_),
    .ZN(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8078_ (.A1(_3160_),
    .A2(_3166_),
    .Z(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8079_ (.A1(_3158_),
    .A2(_3254_),
    .A3(_3255_),
    .ZN(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8080_ (.A1(_3254_),
    .A2(_3256_),
    .ZN(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8081_ (.I(_3236_),
    .ZN(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8082_ (.A1(_3173_),
    .A2(_3258_),
    .ZN(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8083_ (.A1(_3167_),
    .A2(_3237_),
    .B(_3259_),
    .ZN(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8084_ (.A1(_3161_),
    .A2(_3162_),
    .B(_3165_),
    .ZN(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8085_ (.A1(_3184_),
    .A2(_3192_),
    .ZN(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8086_ (.A1(_3184_),
    .A2(_3192_),
    .Z(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8087_ (.A1(_3179_),
    .A2(_3193_),
    .Z(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _8088_ (.A1(_3179_),
    .A2(_3263_),
    .A3(_3264_),
    .B1(_3265_),
    .B2(_3177_),
    .ZN(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8089_ (.A1(_0318_),
    .A2(_1928_),
    .ZN(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8090_ (.A1(_3092_),
    .A2(_3267_),
    .B1(_3183_),
    .B2(_3180_),
    .ZN(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8091_ (.A1(_3266_),
    .A2(_3268_),
    .Z(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8092_ (.A1(_3262_),
    .A2(_3269_),
    .Z(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8093_ (.A1(_3198_),
    .A2(_3235_),
    .ZN(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8094_ (.A1(_3198_),
    .A2(_3235_),
    .ZN(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8095_ (.A1(_3194_),
    .A2(_3272_),
    .B(_3273_),
    .ZN(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8096_ (.A1(_3088_),
    .A2(_3096_),
    .ZN(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8097_ (.A1(_2998_),
    .A2(_3186_),
    .ZN(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8098_ (.A1(_0308_),
    .A2(_1758_),
    .A3(_3275_),
    .B(_3276_),
    .ZN(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8099_ (.A1(_3277_),
    .A2(_3191_),
    .B(_3263_),
    .ZN(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8100_ (.A1(_3203_),
    .A2(_3206_),
    .ZN(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8101_ (.A1(_3203_),
    .A2(_3206_),
    .ZN(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8102_ (.A1(_3201_),
    .A2(_3279_),
    .B(_3280_),
    .ZN(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8103_ (.A1(_0343_),
    .A2(_2099_),
    .ZN(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8104_ (.A1(_0314_),
    .A2(_2011_),
    .ZN(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8105_ (.A1(_3267_),
    .A2(_3284_),
    .ZN(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8106_ (.A1(_3283_),
    .A2(_3285_),
    .Z(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8107_ (.A1(_0577_),
    .A2(_1757_),
    .ZN(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8108_ (.A1(_3186_),
    .A2(_3189_),
    .Z(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8109_ (.A1(_3088_),
    .A2(_3287_),
    .B1(_3288_),
    .B2(_3190_),
    .ZN(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8110_ (.A1(_0443_),
    .A2(_1809_),
    .ZN(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8111_ (.A1(_0409_),
    .A2(_1864_),
    .ZN(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8112_ (.A1(_3287_),
    .A2(_3290_),
    .A3(_3291_),
    .Z(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8113_ (.A1(_3286_),
    .A2(_3289_),
    .A3(_3292_),
    .Z(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8114_ (.A1(_3281_),
    .A2(_3294_),
    .ZN(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8115_ (.A1(_3278_),
    .A2(_3295_),
    .ZN(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8116_ (.A1(_3219_),
    .A2(_3234_),
    .ZN(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8117_ (.A1(_3219_),
    .A2(_3234_),
    .ZN(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8118_ (.A1(_3208_),
    .A2(_3297_),
    .B(_3298_),
    .ZN(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8119_ (.A1(_3225_),
    .A2(_3232_),
    .Z(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8120_ (.A1(_3224_),
    .A2(_3233_),
    .B(_3300_),
    .ZN(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8121_ (.I(_2077_),
    .Z(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8122_ (.A1(_0392_),
    .A2(_3302_),
    .ZN(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8123_ (.A1(_0509_),
    .A2(_1899_),
    .ZN(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8124_ (.A1(_0487_),
    .A2(_1986_),
    .ZN(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8125_ (.A1(_3305_),
    .A2(_3306_),
    .Z(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8126_ (.A1(_3303_),
    .A2(_3307_),
    .Z(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8127_ (.A1(_3228_),
    .A2(_3227_),
    .ZN(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8128_ (.A1(_1371_),
    .A2(\C[0][8] ),
    .A3(_3228_),
    .ZN(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8129_ (.A1(_3309_),
    .A2(_3231_),
    .B(_3310_),
    .ZN(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8130_ (.A1(_0514_),
    .A2(\C[0][9] ),
    .ZN(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8131_ (.A1(_1672_),
    .A2(_3312_),
    .ZN(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8132_ (.A1(_0631_),
    .A2(_1894_),
    .ZN(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8133_ (.I0(_3312_),
    .I1(_3313_),
    .S(_3314_),
    .Z(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8134_ (.A1(_0647_),
    .A2(_1851_),
    .ZN(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8135_ (.A1(_3316_),
    .A2(_3317_),
    .ZN(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8136_ (.A1(_3308_),
    .A2(_3311_),
    .A3(_3318_),
    .Z(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8137_ (.A1(_3301_),
    .A2(_3319_),
    .Z(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8138_ (.A1(_3221_),
    .A2(_3222_),
    .ZN(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8139_ (.A1(_3220_),
    .A2(_3223_),
    .ZN(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8140_ (.A1(_3321_),
    .A2(_3322_),
    .ZN(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8141_ (.A1(_0899_),
    .A2(_2614_),
    .A3(_3128_),
    .ZN(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8142_ (.A1(_3323_),
    .A2(_3324_),
    .Z(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8143_ (.A1(_3320_),
    .A2(_3325_),
    .Z(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _8144_ (.A1(_3296_),
    .A2(_3299_),
    .A3(_3327_),
    .ZN(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8145_ (.A1(_3274_),
    .A2(_3328_),
    .Z(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8146_ (.A1(_3270_),
    .A2(_3329_),
    .Z(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _8147_ (.A1(_3257_),
    .A2(_3261_),
    .A3(_3330_),
    .ZN(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8148_ (.A1(_3253_),
    .A2(_3331_),
    .Z(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8149_ (.A1(_3060_),
    .A2(_3138_),
    .Z(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8150_ (.A1(_3242_),
    .A2(_3333_),
    .B(_3241_),
    .ZN(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8151_ (.A1(_3244_),
    .A2(_3246_),
    .Z(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8152_ (.A1(_3334_),
    .A2(_3335_),
    .Z(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8153_ (.A1(_3332_),
    .A2(_3336_),
    .ZN(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8154_ (.I(_3338_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _8155_ (.A1(_3052_),
    .A2(_3141_),
    .B(_3244_),
    .C(_3140_),
    .ZN(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8156_ (.A1(_3251_),
    .A2(_3252_),
    .B(_3331_),
    .ZN(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8157_ (.A1(_3251_),
    .A2(_3252_),
    .A3(_3331_),
    .ZN(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8158_ (.A1(_3334_),
    .A2(_3340_),
    .B(_3341_),
    .ZN(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8159_ (.A1(_3339_),
    .A2(_3332_),
    .B(_3342_),
    .ZN(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8160_ (.A1(_3261_),
    .A2(_3330_),
    .ZN(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8161_ (.A1(_3261_),
    .A2(_3330_),
    .Z(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8162_ (.A1(_3257_),
    .A2(_3344_),
    .A3(_3345_),
    .ZN(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8163_ (.A1(_3344_),
    .A2(_3346_),
    .ZN(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8164_ (.A1(_3266_),
    .A2(_3268_),
    .ZN(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8165_ (.A1(_3262_),
    .A2(_3269_),
    .ZN(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8166_ (.A1(_3349_),
    .A2(_3350_),
    .ZN(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8167_ (.A1(_3274_),
    .A2(_3328_),
    .ZN(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8168_ (.A1(_3270_),
    .A2(_3329_),
    .ZN(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8169_ (.A1(_3352_),
    .A2(_3353_),
    .ZN(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8170_ (.A1(_3281_),
    .A2(_3294_),
    .ZN(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8171_ (.A1(_3278_),
    .A2(_3295_),
    .B(_3355_),
    .ZN(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _8172_ (.A1(_0897_),
    .A2(_2390_),
    .A3(_3285_),
    .B1(_3284_),
    .B2(_3267_),
    .ZN(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8173_ (.A1(_3356_),
    .A2(_3357_),
    .ZN(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8174_ (.A1(_3299_),
    .A2(_3327_),
    .ZN(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8175_ (.A1(_3299_),
    .A2(_3327_),
    .ZN(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8176_ (.A1(_3296_),
    .A2(_3360_),
    .B(_3361_),
    .ZN(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8177_ (.I(_3289_),
    .ZN(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8178_ (.A1(_3363_),
    .A2(_3292_),
    .ZN(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8179_ (.A1(_3363_),
    .A2(_3292_),
    .ZN(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8180_ (.A1(_3286_),
    .A2(_3364_),
    .B(_3365_),
    .ZN(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8181_ (.A1(_0899_),
    .A2(_2614_),
    .ZN(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _8182_ (.A1(_3204_),
    .A2(_3205_),
    .B1(_3323_),
    .B2(_3367_),
    .ZN(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8183_ (.A1(_0750_),
    .A2(_2101_),
    .ZN(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8184_ (.A1(_3284_),
    .A2(_3370_),
    .ZN(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8185_ (.A1(_0750_),
    .A2(_2013_),
    .B1(_2102_),
    .B2(_0051_),
    .ZN(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8186_ (.A1(_3371_),
    .A2(_3372_),
    .ZN(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8187_ (.A1(_1099_),
    .A2(_1765_),
    .B1(_1810_),
    .B2(_0444_),
    .ZN(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8188_ (.A1(_3992_),
    .A2(_0576_),
    .A3(_3002_),
    .ZN(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8189_ (.A1(_3189_),
    .A2(_3375_),
    .ZN(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8190_ (.A1(_3374_),
    .A2(_3291_),
    .B(_3376_),
    .ZN(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8191_ (.A1(_0443_),
    .A2(_2045_),
    .ZN(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8192_ (.A1(_3375_),
    .A2(_3378_),
    .ZN(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8193_ (.A1(_0408_),
    .A2(_1929_),
    .ZN(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8194_ (.A1(_3379_),
    .A2(_3381_),
    .ZN(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8195_ (.A1(_3377_),
    .A2(_3382_),
    .Z(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8196_ (.A1(_3373_),
    .A2(_3383_),
    .Z(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8197_ (.A1(_3368_),
    .A2(_3384_),
    .Z(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8198_ (.A1(_3366_),
    .A2(_3385_),
    .ZN(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8199_ (.A1(_3301_),
    .A2(_3319_),
    .ZN(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8200_ (.A1(_3320_),
    .A2(_3325_),
    .B(_3387_),
    .ZN(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8201_ (.A1(_0775_),
    .A2(_2562_),
    .A3(_3307_),
    .ZN(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8202_ (.A1(_3305_),
    .A2(_3306_),
    .B(_3389_),
    .ZN(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8203_ (.A1(_3311_),
    .A2(_3318_),
    .ZN(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8204_ (.A1(_3311_),
    .A2(_3318_),
    .ZN(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8205_ (.A1(_3308_),
    .A2(_3392_),
    .B(_3393_),
    .ZN(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8206_ (.A1(_0632_),
    .A2(_1975_),
    .B(_3313_),
    .ZN(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8207_ (.A1(_3312_),
    .A2(_3314_),
    .Z(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8208_ (.A1(_3395_),
    .A2(_3317_),
    .B(_3396_),
    .ZN(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8209_ (.A1(_1178_),
    .A2(\C[0][10] ),
    .ZN(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8210_ (.A1(_1181_),
    .A2(_3398_),
    .ZN(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8211_ (.A1(_0630_),
    .A2(_2275_),
    .ZN(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8212_ (.I0(_3398_),
    .I1(_3399_),
    .S(_3400_),
    .Z(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8213_ (.A1(_0633_),
    .A2(_2250_),
    .ZN(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8214_ (.A1(_3401_),
    .A2(_3403_),
    .ZN(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8215_ (.A1(_3397_),
    .A2(_3404_),
    .Z(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8216_ (.A1(_0390_),
    .A2(_2152_),
    .ZN(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8217_ (.A1(_0720_),
    .A2(_1987_),
    .ZN(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8218_ (.A1(_0488_),
    .A2(_3302_),
    .ZN(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8219_ (.A1(_3407_),
    .A2(_3408_),
    .Z(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8220_ (.A1(_3406_),
    .A2(_3409_),
    .Z(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8221_ (.A1(_3405_),
    .A2(_3410_),
    .Z(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _8222_ (.A1(_3390_),
    .A2(_3394_),
    .A3(_3411_),
    .ZN(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8223_ (.A1(_3388_),
    .A2(_3412_),
    .ZN(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8224_ (.A1(_3386_),
    .A2(_3414_),
    .Z(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8225_ (.A1(_3362_),
    .A2(_3415_),
    .ZN(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8226_ (.A1(_3359_),
    .A2(_3416_),
    .Z(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8227_ (.A1(_3354_),
    .A2(_3417_),
    .Z(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8228_ (.A1(_3351_),
    .A2(_3418_),
    .ZN(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8229_ (.A1(_3348_),
    .A2(_3419_),
    .ZN(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8230_ (.A1(_3343_),
    .A2(_3420_),
    .Z(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8231_ (.I(_3421_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8232_ (.A1(_3344_),
    .A2(_3346_),
    .B(_3419_),
    .ZN(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _8233_ (.A1(_3343_),
    .A2(_3420_),
    .B(_3422_),
    .ZN(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8234_ (.A1(_3354_),
    .A2(_3417_),
    .ZN(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8235_ (.A1(_3351_),
    .A2(_3418_),
    .ZN(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8236_ (.A1(_3425_),
    .A2(_3426_),
    .ZN(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8237_ (.A1(_3356_),
    .A2(_3357_),
    .ZN(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8238_ (.A1(_3362_),
    .A2(_3415_),
    .ZN(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8239_ (.A1(_3359_),
    .A2(_3416_),
    .B(_3429_),
    .ZN(_3430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8240_ (.A1(_3368_),
    .A2(_3384_),
    .ZN(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8241_ (.A1(_3366_),
    .A2(_3385_),
    .ZN(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8242_ (.A1(_3431_),
    .A2(_3432_),
    .ZN(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8243_ (.A1(_3371_),
    .A2(_3433_),
    .ZN(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8244_ (.A1(_3388_),
    .A2(_3412_),
    .ZN(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8245_ (.A1(_3386_),
    .A2(_3414_),
    .ZN(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8246_ (.A1(_3436_),
    .A2(_3437_),
    .ZN(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8247_ (.A1(_3377_),
    .A2(_3382_),
    .ZN(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8248_ (.A1(_3373_),
    .A2(_3383_),
    .ZN(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8249_ (.A1(_3439_),
    .A2(_3440_),
    .ZN(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8250_ (.A1(_1099_),
    .A2(_1949_),
    .ZN(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8251_ (.A1(_0053_),
    .A2(_1931_),
    .A3(_3379_),
    .ZN(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8252_ (.A1(_3290_),
    .A2(_3442_),
    .B(_3443_),
    .ZN(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8253_ (.A1(_0444_),
    .A2(_1930_),
    .ZN(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8254_ (.A1(_3442_),
    .A2(_3446_),
    .ZN(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8255_ (.A1(_0607_),
    .A2(_2123_),
    .ZN(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8256_ (.A1(_3447_),
    .A2(_3448_),
    .Z(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8257_ (.A1(_3444_),
    .A2(_3449_),
    .ZN(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8258_ (.A1(_3370_),
    .A2(_3450_),
    .Z(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8259_ (.A1(_3441_),
    .A2(_3451_),
    .ZN(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8260_ (.A1(_3394_),
    .A2(_3411_),
    .Z(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8261_ (.A1(_3394_),
    .A2(_3411_),
    .Z(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8262_ (.A1(_3390_),
    .A2(_3453_),
    .B(_3454_),
    .ZN(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8263_ (.A1(_3406_),
    .A2(_3409_),
    .ZN(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8264_ (.A1(_3407_),
    .A2(_3408_),
    .B(_3457_),
    .ZN(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8265_ (.A1(_3397_),
    .A2(_3404_),
    .ZN(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8266_ (.A1(_3405_),
    .A2(_3410_),
    .ZN(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8267_ (.A1(_3459_),
    .A2(_3460_),
    .ZN(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8268_ (.I(_0632_),
    .Z(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8269_ (.A1(_3462_),
    .A2(_0003_),
    .B(_3399_),
    .ZN(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8270_ (.A1(_3398_),
    .A2(_3400_),
    .Z(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8271_ (.A1(_3463_),
    .A2(_3403_),
    .B(_3464_),
    .ZN(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8272_ (.A1(_0457_),
    .A2(\C[0][11] ),
    .ZN(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8273_ (.A1(_1672_),
    .A2(_3466_),
    .ZN(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8274_ (.A1(_0631_),
    .A2(_2055_),
    .ZN(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8275_ (.I0(_3466_),
    .I1(_3468_),
    .S(_3469_),
    .Z(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8276_ (.A1(_0718_),
    .A2(_1987_),
    .ZN(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8277_ (.A1(_3470_),
    .A2(_3471_),
    .ZN(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8278_ (.A1(_3465_),
    .A2(_3472_),
    .Z(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8279_ (.A1(_0037_),
    .A2(_3302_),
    .ZN(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8280_ (.A1(_0384_),
    .A2(_2501_),
    .ZN(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8281_ (.A1(_3474_),
    .A2(_3475_),
    .Z(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8282_ (.A1(_3473_),
    .A2(_3476_),
    .Z(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _8283_ (.A1(_3458_),
    .A2(_3461_),
    .A3(_3477_),
    .ZN(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8284_ (.A1(_3455_),
    .A2(_3479_),
    .ZN(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8285_ (.A1(_3438_),
    .A2(_3452_),
    .A3(_3480_),
    .Z(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8286_ (.A1(_3435_),
    .A2(_3481_),
    .Z(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8287_ (.A1(_3430_),
    .A2(_3482_),
    .ZN(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8288_ (.A1(_3428_),
    .A2(_3483_),
    .Z(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8289_ (.A1(_3427_),
    .A2(_3484_),
    .ZN(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8290_ (.A1(_3424_),
    .A2(_3485_),
    .Z(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8291_ (.I(_3486_),
    .Z(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8292_ (.A1(_3371_),
    .A2(_3433_),
    .ZN(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8293_ (.I(_3487_),
    .ZN(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8294_ (.A1(_3452_),
    .A2(_3480_),
    .ZN(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8295_ (.A1(_3452_),
    .A2(_3480_),
    .Z(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _8296_ (.A1(_3438_),
    .A2(_3490_),
    .A3(_3491_),
    .B1(_3481_),
    .B2(_3435_),
    .ZN(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8297_ (.A1(_3441_),
    .A2(_3451_),
    .ZN(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8298_ (.A1(_3455_),
    .A2(_3479_),
    .ZN(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8299_ (.A1(_3494_),
    .A2(_3490_),
    .ZN(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8300_ (.A1(_1094_),
    .A2(_1931_),
    .ZN(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8301_ (.A1(_3378_),
    .A2(_3496_),
    .B1(_3447_),
    .B2(_3448_),
    .ZN(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8302_ (.A1(_0053_),
    .A2(_2203_),
    .ZN(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8303_ (.A1(_0445_),
    .A2(_2579_),
    .Z(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8304_ (.A1(_3496_),
    .A2(_3500_),
    .Z(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8305_ (.A1(_3498_),
    .A2(_3501_),
    .Z(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8306_ (.A1(_3497_),
    .A2(_3502_),
    .ZN(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8307_ (.A1(_3370_),
    .A2(_3450_),
    .ZN(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8308_ (.A1(_3444_),
    .A2(_3449_),
    .B(_3504_),
    .ZN(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8309_ (.A1(_3503_),
    .A2(_3505_),
    .Z(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8310_ (.A1(_3503_),
    .A2(_3505_),
    .ZN(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8311_ (.A1(_3506_),
    .A2(_3507_),
    .ZN(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8312_ (.A1(_3461_),
    .A2(_3477_),
    .Z(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8313_ (.A1(_3461_),
    .A2(_3477_),
    .Z(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8314_ (.A1(_3458_),
    .A2(_3509_),
    .B(_3511_),
    .ZN(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8315_ (.A1(_3474_),
    .A2(_3475_),
    .Z(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8316_ (.A1(_3465_),
    .A2(_3472_),
    .ZN(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8317_ (.A1(_3473_),
    .A2(_3476_),
    .ZN(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8318_ (.A1(_3514_),
    .A2(_3515_),
    .ZN(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8319_ (.A1(_0481_),
    .A2(_2614_),
    .ZN(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8320_ (.I(_0506_),
    .Z(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8321_ (.A1(_3518_),
    .A2(_0005_),
    .A3(_3470_),
    .ZN(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8322_ (.A1(_3466_),
    .A2(_3469_),
    .B(_3519_),
    .ZN(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8323_ (.A1(_0457_),
    .A2(\C[0][12] ),
    .ZN(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8324_ (.A1(_1672_),
    .A2(_3521_),
    .ZN(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8325_ (.A1(_0631_),
    .A2(_2087_),
    .ZN(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8326_ (.I0(_3521_),
    .I1(_3522_),
    .S(_3523_),
    .Z(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8327_ (.A1(_0038_),
    .A2(_3302_),
    .ZN(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8328_ (.A1(_3524_),
    .A2(_3525_),
    .ZN(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8329_ (.A1(_3520_),
    .A2(_3526_),
    .Z(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8330_ (.A1(_3517_),
    .A2(_3527_),
    .ZN(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8331_ (.A1(_3516_),
    .A2(_3528_),
    .ZN(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8332_ (.A1(_3513_),
    .A2(_3529_),
    .ZN(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8333_ (.A1(_3512_),
    .A2(_3530_),
    .ZN(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8334_ (.A1(_3495_),
    .A2(_3508_),
    .A3(_3532_),
    .Z(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8335_ (.A1(_3493_),
    .A2(_3533_),
    .Z(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8336_ (.A1(_3492_),
    .A2(_3534_),
    .Z(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8337_ (.A1(_3489_),
    .A2(_3535_),
    .Z(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8338_ (.A1(_3430_),
    .A2(_3482_),
    .ZN(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8339_ (.A1(_3428_),
    .A2(_3483_),
    .B(_3537_),
    .ZN(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8340_ (.A1(_3536_),
    .A2(_3538_),
    .Z(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8341_ (.A1(_3427_),
    .A2(_3484_),
    .ZN(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8342_ (.A1(_3424_),
    .A2(_3485_),
    .B(_3540_),
    .ZN(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8343_ (.A1(_3539_),
    .A2(_3541_),
    .Z(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8344_ (.I(_3543_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8345_ (.A1(_3492_),
    .A2(_3534_),
    .ZN(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8346_ (.A1(_3489_),
    .A2(_3535_),
    .ZN(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8347_ (.I(_3506_),
    .ZN(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8348_ (.A1(_3512_),
    .A2(_3530_),
    .ZN(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8349_ (.A1(_3508_),
    .A2(_3532_),
    .ZN(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8350_ (.A1(_3547_),
    .A2(_3548_),
    .ZN(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8351_ (.A1(_3520_),
    .A2(_3526_),
    .ZN(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8352_ (.I(_2665_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8353_ (.A1(_0481_),
    .A2(_0007_),
    .A3(_3527_),
    .ZN(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8354_ (.A1(_3550_),
    .A2(_3552_),
    .ZN(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8355_ (.A1(_3518_),
    .A2(_0006_),
    .A3(_3524_),
    .ZN(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8356_ (.A1(_3521_),
    .A2(_3523_),
    .B(_3554_),
    .ZN(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8357_ (.A1(_1528_),
    .A2(\C[0][13] ),
    .ZN(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8358_ (.A1(_1673_),
    .A2(_3556_),
    .ZN(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8359_ (.A1(_3462_),
    .A2(_0006_),
    .ZN(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8360_ (.I0(_3556_),
    .I1(_3557_),
    .S(_3558_),
    .Z(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8361_ (.A1(_3518_),
    .A2(_2665_),
    .ZN(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8362_ (.A1(_3559_),
    .A2(_3560_),
    .ZN(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8363_ (.A1(_3555_),
    .A2(_3561_),
    .Z(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8364_ (.A1(_3553_),
    .A2(_3563_),
    .Z(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8365_ (.A1(_3516_),
    .A2(_3528_),
    .ZN(_3565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8366_ (.A1(_3513_),
    .A2(_3529_),
    .B(_3565_),
    .ZN(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8367_ (.A1(_3564_),
    .A2(_3566_),
    .ZN(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8368_ (.A1(_3497_),
    .A2(_3502_),
    .ZN(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8369_ (.I(_1094_),
    .Z(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8370_ (.A1(_0055_),
    .A2(_0014_),
    .ZN(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8371_ (.A1(_0687_),
    .A2(_2103_),
    .ZN(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _8372_ (.A1(_3446_),
    .A2(_3569_),
    .B1(_3501_),
    .B2(_3498_),
    .ZN(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _8373_ (.A1(_3569_),
    .A2(_3570_),
    .A3(_3571_),
    .ZN(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8374_ (.A1(_3568_),
    .A2(_3573_),
    .ZN(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8375_ (.A1(_3567_),
    .A2(_3574_),
    .ZN(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8376_ (.A1(_3549_),
    .A2(_3575_),
    .Z(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8377_ (.A1(_3546_),
    .A2(_3576_),
    .Z(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8378_ (.A1(_3508_),
    .A2(_3532_),
    .Z(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _8379_ (.A1(_3495_),
    .A2(_3548_),
    .A3(_3578_),
    .B1(_3533_),
    .B2(_3493_),
    .ZN(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8380_ (.A1(_3577_),
    .A2(_3579_),
    .ZN(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _8381_ (.A1(_3544_),
    .A2(_3545_),
    .A3(_3580_),
    .Z(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8382_ (.A1(_3544_),
    .A2(_3545_),
    .B(_3580_),
    .ZN(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8383_ (.A1(_3581_),
    .A2(_3582_),
    .ZN(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8384_ (.A1(_3536_),
    .A2(_3538_),
    .Z(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8385_ (.A1(_3539_),
    .A2(_3541_),
    .B(_3585_),
    .ZN(_3586_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8386_ (.A1(_3584_),
    .A2(_3586_),
    .ZN(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8387_ (.I(_3587_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8388_ (.A1(_3577_),
    .A2(_3579_),
    .ZN(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8389_ (.A1(_3568_),
    .A2(_3573_),
    .ZN(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8390_ (.A1(_3569_),
    .A2(_3570_),
    .ZN(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _8391_ (.A1(_0055_),
    .A2(_0015_),
    .A3(_3500_),
    .ZN(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _8392_ (.A1(_3590_),
    .A2(_3591_),
    .A3(_3571_),
    .ZN(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8393_ (.A1(_0055_),
    .A2(_0015_),
    .ZN(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8394_ (.A1(_3500_),
    .A2(_3594_),
    .ZN(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8395_ (.A1(_3592_),
    .A2(_3595_),
    .Z(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8396_ (.A1(_3518_),
    .A2(_0007_),
    .A3(_3559_),
    .ZN(_3597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8397_ (.A1(_3556_),
    .A2(_3558_),
    .B(_3597_),
    .ZN(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8398_ (.A1(_1597_),
    .A2(\C[0][14] ),
    .ZN(_3599_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8399_ (.A1(_1673_),
    .A2(_3599_),
    .ZN(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8400_ (.A1(_3462_),
    .A2(_2665_),
    .ZN(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8401_ (.I0(_3599_),
    .I1(_3600_),
    .S(_3601_),
    .Z(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8402_ (.A1(_3598_),
    .A2(_3602_),
    .Z(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8403_ (.I(_3603_),
    .ZN(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8404_ (.A1(_3555_),
    .A2(_3561_),
    .ZN(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8405_ (.A1(_3553_),
    .A2(_3563_),
    .ZN(_3607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8406_ (.A1(_3606_),
    .A2(_3607_),
    .ZN(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8407_ (.A1(_3605_),
    .A2(_3608_),
    .Z(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8408_ (.A1(_3596_),
    .A2(_3609_),
    .Z(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8409_ (.A1(_3564_),
    .A2(_3566_),
    .ZN(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8410_ (.A1(_3567_),
    .A2(_3574_),
    .B(_3611_),
    .ZN(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _8411_ (.A1(_3589_),
    .A2(_3610_),
    .A3(_3612_),
    .ZN(_3613_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8412_ (.A1(_3549_),
    .A2(_3575_),
    .ZN(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8413_ (.A1(_3546_),
    .A2(_3576_),
    .B(_3614_),
    .ZN(_3616_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8414_ (.A1(_3613_),
    .A2(_3616_),
    .ZN(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8415_ (.A1(_3588_),
    .A2(_3617_),
    .ZN(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8416_ (.A1(_3539_),
    .A2(_3541_),
    .B(_3582_),
    .C(_3585_),
    .ZN(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8417_ (.A1(_3581_),
    .A2(_3619_),
    .ZN(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8418_ (.A1(_3618_),
    .A2(_3620_),
    .ZN(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8419_ (.I(_3621_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8420_ (.A1(_3588_),
    .A2(_3617_),
    .ZN(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8421_ (.A1(_3581_),
    .A2(_3618_),
    .A3(_3619_),
    .ZN(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8422_ (.A1(_3622_),
    .A2(_3623_),
    .ZN(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8423_ (.A1(_3613_),
    .A2(_3616_),
    .ZN(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8424_ (.A1(_3500_),
    .A2(_3594_),
    .A3(_3592_),
    .ZN(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8425_ (.A1(_3610_),
    .A2(_3612_),
    .Z(_3628_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8426_ (.A1(_3610_),
    .A2(_3612_),
    .Z(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8427_ (.A1(_3589_),
    .A2(_3628_),
    .B(_3629_),
    .ZN(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8428_ (.A1(_3607_),
    .A2(_3605_),
    .B1(_3609_),
    .B2(_3596_),
    .ZN(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8429_ (.A1(_3555_),
    .A2(_3561_),
    .A3(_3603_),
    .ZN(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8430_ (.A1(_3598_),
    .A2(_3602_),
    .ZN(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8431_ (.A1(_3601_),
    .A2(_3599_),
    .B(_3633_),
    .ZN(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8432_ (.A1(\C[0][15] ),
    .A2(_1628_),
    .ZN(_3635_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8433_ (.A1(_3634_),
    .A2(_3635_),
    .Z(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8434_ (.A1(_3632_),
    .A2(_3637_),
    .Z(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8435_ (.A1(_3632_),
    .A2(_3637_),
    .ZN(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8436_ (.A1(_3638_),
    .A2(_3639_),
    .ZN(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8437_ (.A1(_3591_),
    .A2(_3640_),
    .Z(_3641_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8438_ (.A1(_3631_),
    .A2(_3641_),
    .Z(_3642_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8439_ (.A1(_3627_),
    .A2(_3630_),
    .A3(_3642_),
    .Z(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8440_ (.A1(_3626_),
    .A2(_3643_),
    .ZN(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8441_ (.A1(_3624_),
    .A2(_3644_),
    .Z(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8442_ (.I(_3645_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8443_ (.A1(_3626_),
    .A2(_3622_),
    .ZN(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8444_ (.A1(_3643_),
    .A2(_3647_),
    .ZN(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8445_ (.A1(_3623_),
    .A2(_3644_),
    .B(_3648_),
    .ZN(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8446_ (.A1(_3633_),
    .A2(_3635_),
    .B1(_3640_),
    .B2(_3591_),
    .C(_3638_),
    .ZN(_3650_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8447_ (.A1(\C[0][15] ),
    .A2(_3462_),
    .A3(_0007_),
    .A4(_3600_),
    .ZN(_3651_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8448_ (.A1(_1688_),
    .A2(\C[0][16] ),
    .Z(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8449_ (.A1(\C[0][16] ),
    .A2(_1628_),
    .A3(_3651_),
    .ZN(_3653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8450_ (.A1(_3651_),
    .A2(_3652_),
    .B(_3653_),
    .ZN(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8451_ (.A1(_3650_),
    .A2(_3654_),
    .ZN(_3655_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8452_ (.A1(_3627_),
    .A2(_3642_),
    .ZN(_3656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8453_ (.A1(_3627_),
    .A2(_3642_),
    .ZN(_3657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8454_ (.A1(_3631_),
    .A2(_3641_),
    .ZN(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8455_ (.A1(_3630_),
    .A2(_3656_),
    .B(_3657_),
    .C(_3658_),
    .ZN(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _8456_ (.A1(_3649_),
    .A2(_3655_),
    .A3(_3659_),
    .ZN(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8457_ (.I(_3660_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8458_ (.I(_0937_),
    .Z(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8459_ (.A1(_3661_),
    .A2(_3799_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8460_ (.A1(_0937_),
    .A2(_3981_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8461_ (.A1(_3661_),
    .A2(_0181_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8462_ (.A1(_3661_),
    .A2(_3790_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8463_ (.A1(_3661_),
    .A2(_3796_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8464_ (.I(net14),
    .ZN(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8465_ (.I(net13),
    .ZN(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8466_ (.A1(_3663_),
    .A2(_3664_),
    .ZN(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8467_ (.I(_3665_),
    .Z(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8468_ (.I(net13),
    .Z(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8469_ (.A1(_3663_),
    .A2(_3667_),
    .ZN(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8470_ (.I(_3668_),
    .Z(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8471_ (.I(_3668_),
    .Z(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8472_ (.A1(_1696_),
    .A2(_1697_),
    .B(_3670_),
    .ZN(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8473_ (.I(net14),
    .Z(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8474_ (.I(_3664_),
    .Z(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8475_ (.A1(_3673_),
    .A2(_3674_),
    .ZN(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8476_ (.I(_3675_),
    .Z(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8477_ (.A1(_0124_),
    .A2(_3669_),
    .B(_3671_),
    .C(_3676_),
    .ZN(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8478_ (.I(_3667_),
    .Z(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8479_ (.I(_3673_),
    .Z(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8480_ (.A1(_3678_),
    .A2(_0094_),
    .B(_3679_),
    .ZN(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8481_ (.A1(_3660_),
    .A2(_3666_),
    .B1(_3677_),
    .B2(_3680_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8482_ (.I(_3675_),
    .Z(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8483_ (.I(_3663_),
    .Z(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8484_ (.A1(_3683_),
    .A2(_3674_),
    .ZN(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8485_ (.A1(_0066_),
    .A2(_3681_),
    .B1(_3684_),
    .B2(_0064_),
    .ZN(_3685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8486_ (.A1(_3673_),
    .A2(_3667_),
    .ZN(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8487_ (.I(_3686_),
    .Z(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8488_ (.A1(_0068_),
    .A2(_3687_),
    .B1(_3669_),
    .B2(_0070_),
    .ZN(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8489_ (.A1(_3685_),
    .A2(_3688_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8490_ (.A1(_0071_),
    .A2(_3669_),
    .ZN(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _8491_ (.A1(_0069_),
    .A2(_3687_),
    .B1(_3684_),
    .B2(_0065_),
    .C1(_3676_),
    .C2(_0067_),
    .ZN(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8492_ (.A1(_3689_),
    .A2(_3690_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8493_ (.A1(_3683_),
    .A2(_3667_),
    .ZN(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8494_ (.I(_3692_),
    .Z(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8495_ (.A1(_3673_),
    .A2(_3674_),
    .ZN(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8496_ (.I(_3694_),
    .Z(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8497_ (.A1(_0087_),
    .A2(_3693_),
    .B1(_3695_),
    .B2(_0117_),
    .ZN(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8498_ (.A1(_3679_),
    .A2(_3678_),
    .ZN(_3697_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8499_ (.A1(_0102_),
    .A2(_3666_),
    .B1(_3697_),
    .B2(_0072_),
    .ZN(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8500_ (.A1(_3696_),
    .A2(_3698_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8501_ (.I0(_0080_),
    .I1(_0125_),
    .S(_3668_),
    .Z(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8502_ (.A1(_0095_),
    .A2(_3676_),
    .Z(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8503_ (.A1(_3692_),
    .A2(_3699_),
    .B(_3700_),
    .C(_3686_),
    .ZN(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8504_ (.A1(_0110_),
    .A2(_3666_),
    .ZN(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8505_ (.A1(_3702_),
    .A2(_3703_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8506_ (.I(_3674_),
    .Z(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _8507_ (.I0(_0096_),
    .I1(_0111_),
    .I2(_0081_),
    .I3(_0126_),
    .S0(_3704_),
    .S1(_3679_),
    .Z(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8508_ (.I(_3705_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _8509_ (.I0(_0097_),
    .I1(_0112_),
    .I2(_0082_),
    .I3(_0127_),
    .S0(_3704_),
    .S1(_3679_),
    .Z(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8510_ (.I(_3706_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8511_ (.A1(_0098_),
    .A2(_3681_),
    .ZN(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8512_ (.I(_3686_),
    .Z(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _8513_ (.A1(_0113_),
    .A2(_3708_),
    .B1(_3669_),
    .B2(_0128_),
    .C1(_3684_),
    .C2(_0083_),
    .ZN(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8514_ (.A1(_3707_),
    .A2(_3710_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8515_ (.A1(_0084_),
    .A2(_3695_),
    .ZN(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8516_ (.A1(_0129_),
    .A2(_3670_),
    .ZN(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8517_ (.A1(_3692_),
    .A2(_3711_),
    .A3(_3712_),
    .ZN(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8518_ (.I(_3665_),
    .Z(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8519_ (.A1(_0099_),
    .A2(_3693_),
    .B(_3713_),
    .C(_3714_),
    .ZN(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8520_ (.A1(_0114_),
    .A2(_3687_),
    .ZN(_3716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8521_ (.A1(_3715_),
    .A2(_3716_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _8522_ (.I0(_0085_),
    .I1(_0100_),
    .I2(_0130_),
    .I3(_0115_),
    .S0(_3683_),
    .S1(_3704_),
    .Z(_3717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8523_ (.I(_3717_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8524_ (.I(_3683_),
    .Z(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8525_ (.A1(_3719_),
    .A2(_0101_),
    .ZN(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8526_ (.A1(_3675_),
    .A2(_3668_),
    .ZN(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8527_ (.A1(_0131_),
    .A2(_3670_),
    .B1(_3721_),
    .B2(_0086_),
    .ZN(_3722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8528_ (.A1(_3720_),
    .A2(_3722_),
    .ZN(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8529_ (.I0(_0116_),
    .I1(_3723_),
    .S(_3714_),
    .Z(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8530_ (.I(_3724_),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8531_ (.I0(_0118_),
    .I1(_0073_),
    .S(_3694_),
    .Z(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8532_ (.A1(_3692_),
    .A2(_3725_),
    .B(_3708_),
    .ZN(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8533_ (.A1(_0088_),
    .A2(_3681_),
    .ZN(_3728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8534_ (.A1(_0103_),
    .A2(_3666_),
    .ZN(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8535_ (.A1(_3726_),
    .A2(_3728_),
    .B(_3729_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _8536_ (.I0(_0119_),
    .I1(_0074_),
    .I2(_0104_),
    .I3(_0089_),
    .S0(_3678_),
    .S1(_3719_),
    .Z(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8537_ (.I(_3730_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _8538_ (.I0(_0120_),
    .I1(_0075_),
    .I2(_0105_),
    .I3(_0090_),
    .S0(_3678_),
    .S1(_3719_),
    .Z(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8539_ (.I(_3731_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8540_ (.A1(_0091_),
    .A2(_3676_),
    .ZN(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8541_ (.I0(_0121_),
    .I1(_0076_),
    .S(_3695_),
    .Z(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8542_ (.A1(_3693_),
    .A2(_3733_),
    .B(_3708_),
    .ZN(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8543_ (.A1(_0106_),
    .A2(_3714_),
    .ZN(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8544_ (.A1(_3732_),
    .A2(_3734_),
    .B(_3736_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8545_ (.A1(_3719_),
    .A2(_0092_),
    .ZN(_3737_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8546_ (.I0(_0122_),
    .I1(_0077_),
    .S(_3695_),
    .Z(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8547_ (.A1(_3693_),
    .A2(_3738_),
    .B(_3708_),
    .ZN(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8548_ (.A1(_0107_),
    .A2(_3714_),
    .ZN(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8549_ (.A1(_3737_),
    .A2(_3739_),
    .B(_3740_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8550_ (.A1(_1666_),
    .A2(_1667_),
    .B(_3675_),
    .C(_3670_),
    .ZN(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8551_ (.A1(_3704_),
    .A2(_0123_),
    .B(_3686_),
    .C(_3741_),
    .ZN(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8552_ (.A1(_0093_),
    .A2(_3681_),
    .ZN(_3743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8553_ (.A1(_3645_),
    .A2(_3687_),
    .B1(_3742_),
    .B2(_3743_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8554_ (.D(_0132_),
    .CLK(clknet_4_14_0_Clock),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8555_ (.D(_0000_),
    .CLK(clknet_4_2_0_Clock),
    .Q(\A[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8556_ (.D(_0001_),
    .CLK(clknet_4_2_0_Clock),
    .Q(\A[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8557_ (.D(_0002_),
    .CLK(clknet_4_2_0_Clock),
    .Q(\A[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8558_ (.D(_0003_),
    .CLK(clknet_4_8_0_Clock),
    .Q(\A[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8559_ (.D(_0004_),
    .CLK(clknet_4_8_0_Clock),
    .Q(\A[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8560_ (.D(_0005_),
    .CLK(clknet_4_10_0_Clock),
    .Q(\A[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8561_ (.D(_0006_),
    .CLK(clknet_4_10_0_Clock),
    .Q(\A[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8562_ (.D(_0007_),
    .CLK(clknet_4_10_0_Clock),
    .Q(\A[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8563_ (.D(_0008_),
    .CLK(clknet_4_0_0_Clock),
    .Q(\A[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8564_ (.D(_0009_),
    .CLK(clknet_4_1_0_Clock),
    .Q(\A[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8565_ (.D(_0010_),
    .CLK(clknet_4_0_0_Clock),
    .Q(\A[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8566_ (.D(_0011_),
    .CLK(clknet_4_0_0_Clock),
    .Q(\A[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8567_ (.D(_0012_),
    .CLK(clknet_4_0_0_Clock),
    .Q(\A[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8568_ (.D(_0013_),
    .CLK(clknet_4_3_0_Clock),
    .Q(\A[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8569_ (.D(_0014_),
    .CLK(clknet_4_3_0_Clock),
    .Q(\A[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8570_ (.D(_0015_),
    .CLK(clknet_4_3_0_Clock),
    .Q(\A[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8571_ (.D(_0016_),
    .CLK(clknet_4_6_0_Clock),
    .Q(\A[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8572_ (.D(_0017_),
    .CLK(clknet_4_3_0_Clock),
    .Q(\A[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8573_ (.D(_0018_),
    .CLK(clknet_4_3_0_Clock),
    .Q(\A[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8574_ (.D(_0019_),
    .CLK(clknet_4_3_0_Clock),
    .Q(\A[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8575_ (.D(_0020_),
    .CLK(clknet_4_1_0_Clock),
    .Q(\A[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8576_ (.D(_0021_),
    .CLK(clknet_4_1_0_Clock),
    .Q(\A[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8577_ (.D(_0022_),
    .CLK(clknet_4_12_0_Clock),
    .Q(\A[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8578_ (.D(_0023_),
    .CLK(clknet_4_1_0_Clock),
    .Q(\A[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8579_ (.D(_0024_),
    .CLK(clknet_4_6_0_Clock),
    .Q(\A[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8580_ (.D(_0025_),
    .CLK(clknet_4_1_0_Clock),
    .Q(\A[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8581_ (.D(_0026_),
    .CLK(clknet_4_4_0_Clock),
    .Q(\A[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8582_ (.D(_0027_),
    .CLK(clknet_4_4_0_Clock),
    .Q(\A[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8583_ (.D(_0028_),
    .CLK(clknet_4_4_0_Clock),
    .Q(\A[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8584_ (.D(_0029_),
    .CLK(clknet_4_4_0_Clock),
    .Q(\A[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8585_ (.D(_0030_),
    .CLK(clknet_4_6_0_Clock),
    .Q(\A[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8586_ (.D(_0031_),
    .CLK(clknet_4_6_0_Clock),
    .Q(\A[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8587_ (.D(_0032_),
    .CLK(clknet_4_1_0_Clock),
    .Q(\B[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8588_ (.D(_0033_),
    .CLK(clknet_4_2_0_Clock),
    .Q(\B[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8589_ (.D(_0034_),
    .CLK(clknet_4_2_0_Clock),
    .Q(\B[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8590_ (.D(_0035_),
    .CLK(clknet_4_2_0_Clock),
    .Q(\B[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8591_ (.D(_0036_),
    .CLK(clknet_4_9_0_Clock),
    .Q(\B[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8592_ (.D(_0037_),
    .CLK(clknet_4_10_0_Clock),
    .Q(\B[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8593_ (.D(_0038_),
    .CLK(clknet_4_10_0_Clock),
    .Q(\B[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8594_ (.D(_0039_),
    .CLK(clknet_4_10_0_Clock),
    .Q(\B[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8595_ (.D(_0040_),
    .CLK(clknet_4_0_0_Clock),
    .Q(\B[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8596_ (.D(_0041_),
    .CLK(clknet_4_3_0_Clock),
    .Q(\B[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8597_ (.D(_0042_),
    .CLK(clknet_4_3_0_Clock),
    .Q(\B[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8598_ (.D(_0043_),
    .CLK(clknet_4_9_0_Clock),
    .Q(\B[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8599_ (.D(_0044_),
    .CLK(clknet_4_3_0_Clock),
    .Q(\B[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8600_ (.D(_0045_),
    .CLK(clknet_4_9_0_Clock),
    .Q(\B[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8601_ (.D(_0046_),
    .CLK(clknet_4_3_0_Clock),
    .Q(\B[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8602_ (.D(_0047_),
    .CLK(clknet_4_9_0_Clock),
    .Q(\B[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8603_ (.D(_0048_),
    .CLK(clknet_4_0_0_Clock),
    .Q(\B[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8604_ (.D(_0049_),
    .CLK(clknet_4_1_0_Clock),
    .Q(\B[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8605_ (.D(_0050_),
    .CLK(clknet_4_0_0_Clock),
    .Q(\B[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8606_ (.D(_0051_),
    .CLK(clknet_4_1_0_Clock),
    .Q(\B[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8607_ (.D(_0052_),
    .CLK(clknet_4_1_0_Clock),
    .Q(\B[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8608_ (.D(_0053_),
    .CLK(clknet_4_11_0_Clock),
    .Q(\B[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8609_ (.D(_0054_),
    .CLK(clknet_4_11_0_Clock),
    .Q(\B[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8610_ (.D(_0055_),
    .CLK(clknet_4_11_0_Clock),
    .Q(\B[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8611_ (.D(_0056_),
    .CLK(clknet_4_1_0_Clock),
    .Q(\B[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8612_ (.D(_0057_),
    .CLK(clknet_4_2_0_Clock),
    .Q(\B[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8613_ (.D(_0058_),
    .CLK(clknet_4_1_0_Clock),
    .Q(\B[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8614_ (.D(_0059_),
    .CLK(clknet_4_3_0_Clock),
    .Q(\B[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8615_ (.D(_0060_),
    .CLK(clknet_4_1_0_Clock),
    .Q(\B[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8616_ (.D(_0061_),
    .CLK(clknet_4_1_0_Clock),
    .Q(\B[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8617_ (.D(_0062_),
    .CLK(clknet_4_9_0_Clock),
    .Q(\B[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8618_ (.D(_0063_),
    .CLK(clknet_4_7_0_Clock),
    .Q(\B[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8619_ (.D(_0068_),
    .CLK(clknet_4_1_0_Clock),
    .Q(\C[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8620_ (.D(_0069_),
    .CLK(clknet_4_1_0_Clock),
    .Q(\C[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8621_ (.D(_0102_),
    .CLK(clknet_4_1_0_Clock),
    .Q(\C[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8622_ (.D(_0110_),
    .CLK(clknet_4_1_0_Clock),
    .Q(\C[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8623_ (.D(_0111_),
    .CLK(clknet_4_0_0_Clock),
    .Q(\C[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8624_ (.D(_0112_),
    .CLK(clknet_4_0_0_Clock),
    .Q(\C[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8625_ (.D(_0113_),
    .CLK(clknet_4_2_0_Clock),
    .Q(\C[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8626_ (.D(_0114_),
    .CLK(clknet_4_2_0_Clock),
    .Q(\C[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8627_ (.D(_0115_),
    .CLK(clknet_4_8_0_Clock),
    .Q(\C[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8628_ (.D(_0116_),
    .CLK(clknet_4_8_0_Clock),
    .Q(\C[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8629_ (.D(_0103_),
    .CLK(clknet_4_8_0_Clock),
    .Q(\C[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8630_ (.D(_0104_),
    .CLK(clknet_4_10_0_Clock),
    .Q(\C[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8631_ (.D(_0105_),
    .CLK(clknet_4_10_0_Clock),
    .Q(\C[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8632_ (.D(_0106_),
    .CLK(clknet_4_11_0_Clock),
    .Q(\C[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8633_ (.D(_0107_),
    .CLK(clknet_4_11_0_Clock),
    .Q(\C[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8634_ (.D(_0108_),
    .CLK(clknet_4_11_0_Clock),
    .Q(\C[0][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8635_ (.D(_0109_),
    .CLK(clknet_4_11_0_Clock),
    .Q(\C[0][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8636_ (.D(_0066_),
    .CLK(clknet_4_1_0_Clock),
    .Q(\C[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8637_ (.D(_0067_),
    .CLK(clknet_4_0_0_Clock),
    .Q(\C[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8638_ (.D(_0087_),
    .CLK(clknet_4_9_0_Clock),
    .Q(\C[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8639_ (.D(_0095_),
    .CLK(clknet_4_2_0_Clock),
    .Q(\C[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8640_ (.D(_0096_),
    .CLK(clknet_4_0_0_Clock),
    .Q(\C[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8641_ (.D(_0097_),
    .CLK(clknet_4_0_0_Clock),
    .Q(\C[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8642_ (.D(_0098_),
    .CLK(clknet_4_0_0_Clock),
    .Q(\C[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8643_ (.D(_0099_),
    .CLK(clknet_4_8_0_Clock),
    .Q(\C[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8644_ (.D(_0100_),
    .CLK(clknet_4_8_0_Clock),
    .Q(\C[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8645_ (.D(_0101_),
    .CLK(clknet_4_9_0_Clock),
    .Q(\C[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8646_ (.D(_0088_),
    .CLK(clknet_4_8_0_Clock),
    .Q(\C[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8647_ (.D(_0089_),
    .CLK(clknet_4_10_0_Clock),
    .Q(\C[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8648_ (.D(_0090_),
    .CLK(clknet_4_11_0_Clock),
    .Q(\C[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8649_ (.D(_0091_),
    .CLK(clknet_4_11_0_Clock),
    .Q(\C[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8650_ (.D(_0092_),
    .CLK(clknet_4_11_0_Clock),
    .Q(\C[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8651_ (.D(_0093_),
    .CLK(clknet_4_11_0_Clock),
    .Q(\C[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8652_ (.D(_0094_),
    .CLK(clknet_4_11_0_Clock),
    .Q(\C[1][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8653_ (.D(_0070_),
    .CLK(clknet_4_4_0_Clock),
    .Q(\C[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8654_ (.D(_0071_),
    .CLK(clknet_4_4_0_Clock),
    .Q(\C[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8655_ (.D(_0117_),
    .CLK(clknet_4_12_0_Clock),
    .Q(\C[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8656_ (.D(_0125_),
    .CLK(clknet_4_6_0_Clock),
    .Q(\C[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8657_ (.D(_0126_),
    .CLK(clknet_4_6_0_Clock),
    .Q(\C[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8658_ (.D(_0127_),
    .CLK(clknet_4_6_0_Clock),
    .Q(\C[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8659_ (.D(_0128_),
    .CLK(clknet_4_7_0_Clock),
    .Q(\C[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8660_ (.D(_0129_),
    .CLK(clknet_4_14_0_Clock),
    .Q(\C[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8661_ (.D(_0130_),
    .CLK(clknet_4_12_0_Clock),
    .Q(\C[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8662_ (.D(_0131_),
    .CLK(clknet_4_14_0_Clock),
    .Q(\C[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8663_ (.D(_0118_),
    .CLK(clknet_4_14_0_Clock),
    .Q(\C[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8664_ (.D(_0119_),
    .CLK(clknet_4_15_0_Clock),
    .Q(\C[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8665_ (.D(_0120_),
    .CLK(clknet_4_15_0_Clock),
    .Q(\C[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8666_ (.D(_0121_),
    .CLK(clknet_4_15_0_Clock),
    .Q(\C[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8667_ (.D(_0122_),
    .CLK(clknet_4_15_0_Clock),
    .Q(\C[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8668_ (.D(_0123_),
    .CLK(clknet_4_15_0_Clock),
    .Q(\C[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8669_ (.D(_0124_),
    .CLK(clknet_4_15_0_Clock),
    .Q(\C[2][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8670_ (.D(_0064_),
    .CLK(clknet_4_4_0_Clock),
    .Q(\C[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8671_ (.D(_0065_),
    .CLK(clknet_4_4_0_Clock),
    .Q(\C[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8672_ (.D(_0072_),
    .CLK(clknet_4_4_0_Clock),
    .Q(\C[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8673_ (.D(_0080_),
    .CLK(clknet_4_4_0_Clock),
    .Q(\C[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8674_ (.D(_0081_),
    .CLK(clknet_4_4_0_Clock),
    .Q(\C[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8675_ (.D(_0082_),
    .CLK(clknet_4_5_0_Clock),
    .Q(\C[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8676_ (.D(_0083_),
    .CLK(clknet_4_4_0_Clock),
    .Q(\C[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8677_ (.D(_0084_),
    .CLK(clknet_4_12_0_Clock),
    .Q(\C[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8678_ (.D(_0085_),
    .CLK(clknet_4_7_0_Clock),
    .Q(\C[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8679_ (.D(_0086_),
    .CLK(clknet_4_7_0_Clock),
    .Q(\C[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8680_ (.D(_0073_),
    .CLK(clknet_4_7_0_Clock),
    .Q(\C[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8681_ (.D(_0074_),
    .CLK(clknet_4_7_0_Clock),
    .Q(\C[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8682_ (.D(_0075_),
    .CLK(clknet_4_11_0_Clock),
    .Q(\C[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8683_ (.D(_0076_),
    .CLK(clknet_4_12_0_Clock),
    .Q(\C[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8684_ (.D(_0077_),
    .CLK(clknet_4_12_0_Clock),
    .Q(\C[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8685_ (.D(_0078_),
    .CLK(clknet_4_13_0_Clock),
    .Q(\C[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8686_ (.D(_0079_),
    .CLK(clknet_4_13_0_Clock),
    .Q(\C[3][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8687_ (.D(_0133_),
    .CLK(clknet_4_5_0_Clock),
    .Q(net16));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8688_ (.D(_0134_),
    .CLK(clknet_4_5_0_Clock),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8689_ (.D(_0135_),
    .CLK(clknet_4_5_0_Clock),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8690_ (.D(_0136_),
    .CLK(clknet_4_5_0_Clock),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8691_ (.D(_0137_),
    .CLK(clknet_4_5_0_Clock),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8692_ (.D(_0138_),
    .CLK(clknet_4_5_0_Clock),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8693_ (.D(_0139_),
    .CLK(clknet_4_5_0_Clock),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8694_ (.D(_0140_),
    .CLK(clknet_4_7_0_Clock),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8695_ (.D(_0141_),
    .CLK(clknet_4_7_0_Clock),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8696_ (.D(_0142_),
    .CLK(clknet_4_13_0_Clock),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8697_ (.D(_0143_),
    .CLK(clknet_4_7_0_Clock),
    .Q(net17));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8698_ (.D(_0144_),
    .CLK(clknet_4_12_0_Clock),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8699_ (.D(_0145_),
    .CLK(clknet_4_13_0_Clock),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8700_ (.D(_0146_),
    .CLK(clknet_4_13_0_Clock),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8701_ (.D(_0147_),
    .CLK(clknet_4_13_0_Clock),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _8702_ (.D(_0148_),
    .CLK(clknet_4_13_0_Clock),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_Clock (.I(Clock),
    .Z(clknet_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input1 (.I(Enable),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input2 (.I(K[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input3 (.I(K[1]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input4 (.I(K[2]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(X[0]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(X[1]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(X[2]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(X[3]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(X[4]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(X[5]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(X[6]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input12 (.I(X[7]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(Z[0]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(Z[1]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(reset),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output16 (.I(net16),
    .Z(Result[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output17 (.I(net17),
    .Z(Result[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output18 (.I(net18),
    .Z(Result[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output19 (.I(net19),
    .Z(Result[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output20 (.I(net20),
    .Z(Result[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output21 (.I(net21),
    .Z(Result[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output22 (.I(net22),
    .Z(Result[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output23 (.I(net23),
    .Z(Result[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output24 (.I(net24),
    .Z(Result[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output25 (.I(net25),
    .Z(Result[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output26 (.I(net26),
    .Z(Result[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output27 (.I(net27),
    .Z(Result[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output28 (.I(net28),
    .Z(Result[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output29 (.I(net29),
    .Z(Result[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output30 (.I(net30),
    .Z(Result[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output31 (.I(net31),
    .Z(Result[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output32 (.I(net32),
    .Z(Result[9]));
 gf180mcu_fd_sc_mcu7t5v0__tieh multiply_komal_33 (.Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_Clock (.I(clknet_0_Clock),
    .Z(clknet_3_0_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_Clock (.I(clknet_0_Clock),
    .Z(clknet_3_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_Clock (.I(clknet_0_Clock),
    .Z(clknet_3_2_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_Clock (.I(clknet_0_Clock),
    .Z(clknet_3_3_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_Clock (.I(clknet_0_Clock),
    .Z(clknet_3_4_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_Clock (.I(clknet_0_Clock),
    .Z(clknet_3_5_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_Clock (.I(clknet_0_Clock),
    .Z(clknet_3_6_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_Clock (.I(clknet_0_Clock),
    .Z(clknet_3_7_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_0_0_Clock (.I(clknet_3_0_0_Clock),
    .Z(clknet_4_0_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_1_0_Clock (.I(clknet_3_0_0_Clock),
    .Z(clknet_4_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_2_0_Clock (.I(clknet_3_1_0_Clock),
    .Z(clknet_4_2_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_3_0_Clock (.I(clknet_3_1_0_Clock),
    .Z(clknet_4_3_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_4_0_Clock (.I(clknet_3_2_0_Clock),
    .Z(clknet_4_4_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_5_0_Clock (.I(clknet_3_2_0_Clock),
    .Z(clknet_4_5_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_6_0_Clock (.I(clknet_3_3_0_Clock),
    .Z(clknet_4_6_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_7_0_Clock (.I(clknet_3_3_0_Clock),
    .Z(clknet_4_7_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_8_0_Clock (.I(clknet_3_4_0_Clock),
    .Z(clknet_4_8_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_9_0_Clock (.I(clknet_3_4_0_Clock),
    .Z(clknet_4_9_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_10_0_Clock (.I(clknet_3_5_0_Clock),
    .Z(clknet_4_10_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_11_0_Clock (.I(clknet_3_5_0_Clock),
    .Z(clknet_4_11_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_12_0_Clock (.I(clknet_3_6_0_Clock),
    .Z(clknet_4_12_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_13_0_Clock (.I(clknet_3_6_0_Clock),
    .Z(clknet_4_13_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_14_0_Clock (.I(clknet_3_7_0_Clock),
    .Z(clknet_4_14_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_15_0_Clock (.I(clknet_3_7_0_Clock),
    .Z(clknet_4_15_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer1 (.I(_1790_),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 rebuffer2 (.I(_1874_),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer3 (.I(_1821_),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer4 (.I(net41),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer5 (.I(_1780_),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer6 (.I(_1889_),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlya_1 rebuffer7 (.I(_2189_),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer8 (.I(net42),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 rebuffer9 (.I(_3604_),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer10 (.I(_1713_),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlya_2 rebuffer11 (.I(_3572_),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 rebuffer12 (.I(_0311_),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__B (.I(\A[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6870__I (.I(\A[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__B (.I(\A[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__B (.I(\A[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__B (.I(\A[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7029__B (.I(\A[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__B2 (.I(\A[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__B2 (.I(\A[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__B2 (.I(\A[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__B2 (.I(\A[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__A1 (.I(\A[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__A1 (.I(\A[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__I (.I(\A[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__B2 (.I(\A[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__I (.I(\A[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A1 (.I(\A[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__I (.I(\A[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A3 (.I(\A[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A1 (.I(\A[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__I (.I(\A[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__A1 (.I(\A[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__I (.I(\A[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__B (.I(\A[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__B (.I(\A[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__B (.I(\A[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__B (.I(\A[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__B (.I(\A[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__B (.I(\A[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__B (.I(\A[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__I (.I(\B[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__B2 (.I(\B[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__B (.I(\B[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__B (.I(\B[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__B (.I(\B[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__B (.I(\B[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__B (.I(\B[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A1 (.I(\B[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A1 (.I(\B[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6585__I (.I(\B[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__A1 (.I(\B[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__I (.I(\B[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__A1 (.I(\B[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__I (.I(\B[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A1 (.I(\B[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__I (.I(\B[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__I (.I(\B[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A1 (.I(\B[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__I (.I(\B[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A1 (.I(\B[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__I (.I(\B[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A1 (.I(\B[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__I (.I(\B[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__A3 (.I(\B[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__A1 (.I(\B[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__I (.I(\B[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__B2 (.I(\B[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__B2 (.I(\B[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__B2 (.I(\B[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A3 (.I(\B[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A3 (.I(\B[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A3 (.I(\B[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__B2 (.I(\B[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__B2 (.I(\B[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__A1 (.I(\B[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__B2 (.I(\B[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__B2 (.I(\B[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A1 (.I(\B[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7580__A2 (.I(\C[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__A2 (.I(\C[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__A1 (.I(\C[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7727__A1 (.I(\C[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7857__A2 (.I(\C[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7855__A2 (.I(\C[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7942__I (.I(\C[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8128__A2 (.I(\C[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8050__A2 (.I(\C[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__A2 (.I(\C[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__A2 (.I(\C[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__A2 (.I(\C[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__A2 (.I(\C[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7358__A2 (.I(\C[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__A2 (.I(\C[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__A2 (.I(\C[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__A2 (.I(\C[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__A2 (.I(\C[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6710__A2 (.I(\C[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6775__A2 (.I(\C[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__A2 (.I(\C[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__A2 (.I(\C[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A2 (.I(\C[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__A2 (.I(\C[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A2 (.I(\C[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A2 (.I(\C[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A2 (.I(\C[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__A2 (.I(\C[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__A1 (.I(\C[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A2 (.I(\C[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A1 (.I(\C[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A1 (.I(\C[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A2 (.I(\C[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__A2 (.I(\C[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__A2 (.I(\C[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__A2 (.I(\C[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A1 (.I(\C[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__A1 (.I(\C[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__A1 (.I(\C[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__A2 (.I(\C[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A2 (.I(\C[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A2 (.I(\C[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__A2 (.I(\C[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__A2 (.I(\C[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A2 (.I(\C[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A1 (.I(\C[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__A1 (.I(\C[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A1 (.I(\C[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A1 (.I(\C[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A1 (.I(\C[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A1 (.I(\C[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A2 (.I(\C[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A3 (.I(\C[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__A2 (.I(\C[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A2 (.I(\C[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__A2 (.I(\C[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__A2 (.I(\C[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_Clock_I (.I(Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(Enable));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(K[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(K[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(K[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(X[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(X[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(X[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(X[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(X[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(X[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(X[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(X[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(Z[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(Z[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8555__D (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__A4 (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__A4 (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6592__A2 (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__D (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7713__A2 (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6761__A2 (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__A2 (.I(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8557__D (.I(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7714__A4 (.I(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7713__B1 (.I(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__A2 (.I(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8558__D (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8269__A2 (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7668__A2 (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7224__A2 (.I(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__D (.I(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__A3 (.I(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__B1 (.I(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__A2 (.I(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8560__D (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8321__A2 (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7408__A2 (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__A2 (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__D (.I(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8359__A2 (.I(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8355__A2 (.I(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__A2 (.I(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8562__D (.I(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8447__A3 (.I(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8396__A2 (.I(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8353__A2 (.I(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__D (.I(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__A2 (.I(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__A2 (.I(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__A2 (.I(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8564__D (.I(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7597__A2 (.I(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6682__A2 (.I(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6629__A2 (.I(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__D (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7612__A3 (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__A2 (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__A2 (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8566__D (.I(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7694__A2 (.I(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7646__A2 (.I(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__A3 (.I(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8567__D (.I(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__A2 (.I(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__A2 (.I(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__A2 (.I(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8568__D (.I(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__A2 (.I(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__A2 (.I(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__A2 (.I(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8569__D (.I(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8370__A2 (.I(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__A2 (.I(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__A2 (.I(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8570__D (.I(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8393__A2 (.I(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8391__A2 (.I(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7183__A2 (.I(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8571__D (.I(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__A1 (.I(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A1 (.I(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A1 (.I(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8575__D (.I(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A2 (.I(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__A1 (.I(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A2 (.I(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__D (.I(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__A1 (.I(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__A1 (.I(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A1 (.I(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8577__D (.I(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A1 (.I(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__I (.I(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__D (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__A2 (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__A2 (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A1 (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8579__D (.I(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__A1 (.I(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A1 (.I(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__A1 (.I(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__D (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A1 (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__I (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A1 (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8581__D (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__A1 (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__B2 (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__A1 (.I(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8582__D (.I(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A1 (.I(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A1 (.I(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A1 (.I(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8583__D (.I(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__A1 (.I(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A1 (.I(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A1 (.I(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__D (.I(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__A1 (.I(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__A2 (.I(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A2 (.I(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__D (.I(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A1 (.I(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A2 (.I(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__A2 (.I(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8586__D (.I(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A1 (.I(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A1 (.I(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A1 (.I(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8587__D (.I(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__A2 (.I(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__D (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__A1 (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__A2 (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A2 (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8589__D (.I(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7714__A1 (.I(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A4 (.I(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__B1 (.I(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8590__D (.I(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7724__A1 (.I(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7673__A1 (.I(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__A1 (.I(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8591__D (.I(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A2 (.I(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A4 (.I(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__B1 (.I(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__D (.I(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__A1 (.I(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A2 (.I(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A2 (.I(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8593__D (.I(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8327__A1 (.I(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A2 (.I(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__A2 (.I(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8594__D (.I(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A2 (.I(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A2 (.I(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A2 (.I(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8595__D (.I(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6600__A1 (.I(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__A3 (.I(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__A1 (.I(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8597__D (.I(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__A1 (.I(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__A1 (.I(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A2 (.I(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8598__D (.I(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__A1 (.I(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A1 (.I(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__A1 (.I(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8599__D (.I(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__A1 (.I(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8600__D (.I(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__A1 (.I(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__A1 (.I(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__A2 (.I(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8601__D (.I(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8602__D (.I(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A4 (.I(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8603__D (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7597__A1 (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__A1 (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__A2 (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8604__D (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7994__A1 (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__A1 (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A2 (.I(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8605__D (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__A1 (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7658__A1 (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__A2 (.I(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8606__D (.I(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8185__B2 (.I(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__A2 (.I(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__A2 (.I(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8607__D (.I(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7991__A1 (.I(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__B1 (.I(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A2 (.I(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8608__D (.I(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8302__A1 (.I(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8251__A1 (.I(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A2 (.I(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8609__D (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A2 (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__A1 (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A2 (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8611__D (.I(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A2 (.I(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__A1 (.I(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__A1 (.I(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8612__D (.I(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__A1 (.I(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A2 (.I(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__A2 (.I(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8613__D (.I(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__A1 (.I(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A1 (.I(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A1 (.I(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8614__D (.I(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__B2 (.I(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__A1 (.I(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A1 (.I(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8615__D (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__A1 (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A1 (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A1 (.I(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8616__D (.I(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7425__A1 (.I(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__A1 (.I(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A2 (.I(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8617__D (.I(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7434__A1 (.I(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__A1 (.I(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__A1 (.I(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8618__D (.I(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A2 (.I(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__A2 (.I(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__B2 (.I(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8670__D (.I(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8485__B2 (.I(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8671__D (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__B2 (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8636__D (.I(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8485__A1 (.I(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8637__D (.I(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__C2 (.I(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8619__D (.I(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__A1 (.I(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8620__D (.I(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__A1 (.I(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8653__D (.I(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__B2 (.I(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8672__D (.I(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__B2 (.I(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8680__D (.I(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8531__I1 (.I(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8681__D (.I(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8536__I1 (.I(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8682__D (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8538__I1 (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8683__D (.I(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8541__I1 (.I(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8684__D (.I(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__I1 (.I(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8673__D (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__I0 (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8674__D (.I(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__I2 (.I(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8675__D (.I(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8509__I2 (.I(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8676__D (.I(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__C2 (.I(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8677__D (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8515__A1 (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8678__D (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8522__I0 (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8679__D (.I(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8527__B2 (.I(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8638__D (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8497__A1 (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8646__D (.I(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8533__A1 (.I(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8647__D (.I(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8536__I3 (.I(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8648__D (.I(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8538__I3 (.I(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8649__D (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8540__A1 (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8650__D (.I(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8545__A2 (.I(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8651__D (.I(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8552__A1 (.I(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8652__D (.I(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__A2 (.I(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8639__D (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8502__A1 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8640__D (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__I0 (.I(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8641__D (.I(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8509__I0 (.I(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8642__D (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8511__A1 (.I(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8643__D (.I(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8519__A1 (.I(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8644__D (.I(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8522__I1 (.I(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8645__D (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8525__A2 (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8621__D (.I(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__A1 (.I(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8629__D (.I(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8534__A1 (.I(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8630__D (.I(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8536__I2 (.I(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8631__D (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8538__I2 (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8632__D (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8543__A1 (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8633__D (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8548__A1 (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8622__D (.I(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8504__A1 (.I(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8623__D (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__I1 (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8624__D (.I(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8509__I1 (.I(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8625__D (.I(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__A1 (.I(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8626__D (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8520__A1 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8627__D (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8522__I3 (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8628__D (.I(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8529__I0 (.I(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8655__D (.I(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8497__B2 (.I(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8663__D (.I(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8531__I0 (.I(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8665__D (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8538__I0 (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8666__D (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8541__I0 (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8667__D (.I(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__I0 (.I(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8668__D (.I(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8551__A2 (.I(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8669__D (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8477__A1 (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8657__D (.I(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__I3 (.I(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8658__D (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8509__I3 (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8659__D (.I(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__B2 (.I(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8660__D (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8516__A1 (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8661__D (.I(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8522__I2 (.I(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8662__D (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8527__A1 (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8687__D (.I(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8688__D (.I(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8689__D (.I(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8691__D (.I(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8693__D (.I(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8694__D (.I(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8697__D (.I(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8699__D (.I(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8700__D (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8702__D (.I(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A2 (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__A2 (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__A2 (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__A2 (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__A2 (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__A2 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__A1 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__A1 (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__A2 (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__A1 (.I(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__A2 (.I(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__A1 (.I(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A2 (.I(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8461__A2 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A2 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A2 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__B2 (.I(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__B (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7625__A2 (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7593__A2 (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A2 (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__I (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7477__A3 (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7475__A2 (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__A2 (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__I (.I(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7516__A2 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__I (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__A2 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A2 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__A1 (.I(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__A1 (.I(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A1 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__A1 (.I(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__A2 (.I(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__A1 (.I(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__I (.I(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A1 (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__A1 (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A2 (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__I (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A1 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__A1 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A1 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__I (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__A1 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__A1 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__A1 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A2 (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__A1 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A2 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__I (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A1 (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__A1 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A1 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__A2 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__A1 (.I(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6628__A1 (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A1 (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A2 (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__A2 (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7585__A1 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A1 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A4 (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__A1 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6629__A1 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6604__A1 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A2 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__A1 (.I(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A1 (.I(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7183__A1 (.I(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__I (.I(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__B1 (.I(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__A2 (.I(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A2 (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__I (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__A2 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A2 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A2 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A2 (.I(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6036__A3 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__A2 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__I (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__I (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__A2 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A2 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__A2 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__A2 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__I (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__I (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__B1 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__B1 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__B1 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__B1 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7928__A2 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7838__A2 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__I (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__I (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8098__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8017__A2 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A2 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__A1 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__A1 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A1 (.I(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A1 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__A1 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__I (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A1 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__A1 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7925__A1 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__I (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__I (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A2 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__I (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A2 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A2 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7904__A2 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7822__A2 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__I (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__I (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8009__A1 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A2 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A2 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__I (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A1 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8016__A2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__A2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__I (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__I (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8014__A2 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7837__A1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__A2 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__I (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__A1 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__A1 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A3 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A3 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A3 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__I (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__I (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A3 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__A2 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__A3 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A3 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7623__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__I (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7721__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__I (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__B2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7710__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__I (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__I (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__A3 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__A2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A2 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__B3 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A1 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5671__A1 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A1 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A1 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__I (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__I (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7840__A1 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__I (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__I (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__I (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__A3 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A2 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__A3 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__A3 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__A3 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A3 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7718__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7662__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__A2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7718__A2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7662__A2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__A2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__A2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__A2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__I (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__A4 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__B1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__A4 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__B1 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__B2 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__I (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__A1 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__I (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__A1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__I (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__A2 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A2 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__A3 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__A2 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__I (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__I (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__I (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7924__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__I (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A2 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__A3 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A2 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__A3 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A1 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A1 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A1 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__A1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A2 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__A1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7645__A1 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__A1 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7596__A1 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__I (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A2 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__I (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__I (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__I (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__A2 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A3 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__I (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A3 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A3 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__A2 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__A2 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7852__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7787__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A3 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__A3 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__A3 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A3 (.I(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7852__A2 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7787__A2 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A2 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A2 (.I(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7938__B2 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__A1 (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__I (.I(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__B2 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7792__A1 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A2 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__I (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8280__A1 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8028__A1 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A4 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__B1 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__A1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__B2 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7954__A1 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7793__A1 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__I (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A2 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8216__A1 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A2 (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__I (.I(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7780__A1 (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__I (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__I (.I(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__I (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__A3 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__A1 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__A1 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__I (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__A1 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A1 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__A1 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7780__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__I (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__I (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__A1 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A2 (.I(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8044__A1 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7670__I (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8193__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__I (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__A2 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__I (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8111__A1 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__A2 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8008__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__A3 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A2 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__I (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A3 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__A2 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A3 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__A2 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__A4 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__B1 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__A2 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__I (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__A1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__A2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__A1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__A1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__A1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__B2 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__I (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A2 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__A2 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A2 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__A3 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__B1 (.I(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7959__A1 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__I (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7668__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__I (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7591__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__I (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__B2 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__A1 (.I(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__A1 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8253__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__B2 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__I (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__I (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__A1 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5412__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A3 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__A1 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8050__A1 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__A1 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__I (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__I (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8323__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__A1 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__B2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__I (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__I (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__I (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__I (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A2 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__I (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__A4 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A3 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__B (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A1 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__A3 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__B1 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A3 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A3 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__B1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__A2 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__I (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7608__I (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__I (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__A3 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__B2 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__B2 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__I (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__A3 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A3 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__B2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__B2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7857__A1 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__A1 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__A1 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__A1 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__A3 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__B1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A3 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__A3 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__B2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__I (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__B2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7851__A1 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__A1 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__A1 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7851__A2 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__A2 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__A2 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8353__A1 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8319__A1 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7938__A1 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__A2 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__A2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A3 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__A1 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8046__A1 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A2 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__I (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8218__A1 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7725__A1 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__A2 (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__I (.I(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__A1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__A1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A1 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__B2 (.I(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__I (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A2 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__A2 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__A2 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__A2 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__A2 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__A2 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__A2 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5671__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__A2 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7856__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8320__I (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__A2 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__I (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__I (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8123__A1 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__A2 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__I (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A2 (.I(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__A1 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__A2 (.I(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__A1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__A1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__A1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6710__A1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__A1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__I (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8130__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7855__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8010__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A2 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__A2 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__A2 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__A2 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A4 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__A4 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__B1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__A1 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__A1 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__A2 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A3 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7620__A1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__B1 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__A2 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__A2 (.I(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A1 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__A1 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A2 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A1 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__A3 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__A1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__A2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__A2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__A2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7945__B1 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__A2 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__I (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__I (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__I (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7855__A3 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7791__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__I (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__A2 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__A2 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__I (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__A2 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__A2 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A1 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A1 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__A1 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8188__A2 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8013__A2 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__I (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__I (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8107__A1 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8014__B2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7929__A1 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__A2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A2 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__A2 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__A1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A1 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A1 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A1 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__B (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A1 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A1 (.I(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8255__A1 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__I (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__A2 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A2 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__A1 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A2 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A2 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__A1 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__A1 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8211__A1 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__I (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8268__I (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8206__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__A3 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__A2 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8213__A1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__A1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__A4 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__B1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__A2 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__A1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__A1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__A2 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8134__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A3 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A2 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A3 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__I (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__I (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__I (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A4 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__B1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__I (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__I (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A2 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__A2 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A4 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__B1 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__A3 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__B1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__A3 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__B (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8371__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__I (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5910__A1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A2 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__A1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__A1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A2 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A2 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A2 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A2 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__A1 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8036__A1 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__I (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8276__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8038__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__I (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8217__A1 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__A1 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A2 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__A2 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A2 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A3 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__A2 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A3 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__A2 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__A2 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A3 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__A3 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A3 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8185__A1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8183__A1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__I (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7842__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7708__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__I (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__A2 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__A1 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7657__A1 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__A2 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__A1 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A1 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A3 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__I (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__A3 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5695__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__A2 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__A2 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__B2 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__A2 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7709__A1 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__A2 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A2 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A3 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__A2 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A1 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A1 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__I (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__B2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7726__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__B1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A4 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__A1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__A1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A1 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__A1 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__A2 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A2 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A2 (.I(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__A1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__B (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8030__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7957__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7868__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__I (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__I (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A4 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__B1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A3 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__A2 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__A2 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A2 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7824__A1 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7759__A1 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__A2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__B (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__A1 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__A1 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A1 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__A1 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A3 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__A1 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A1 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A3 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__B (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A3 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__A1 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__A1 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__I (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A3 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__A1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A3 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A2 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__A2 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A2 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__A2 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A2 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__I (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__A3 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__A1 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7770__A1 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7710__A2 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__B2 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__I (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8172__A1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__A1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__A1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5726__A2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8181__A1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8141__A1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7713__A1 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A2 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__I (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7907__A1 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7696__A1 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__I (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A1 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__A1 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A1 (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__A1 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A1 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__A1 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A2 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7581__A1 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A3 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A3 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__A3 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A3 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__A1 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8031__A1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7869__A1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7667__A1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__I (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7714__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7713__B2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__A2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__A2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A3 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8460__A1 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8458__I (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A1 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A1 (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7638__A1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__A1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7551__A2 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__A2 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__I (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A2 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__A2 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A2 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7978__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__A2 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__A2 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5822__A1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__A2 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7277__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__I (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A4 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A2 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A2 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A1 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__A1 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__A2 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5820__A3 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__B (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5976__A2 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__A2 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__A1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__A1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A1 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A2 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A1 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A3 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A1 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__A1 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7299__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7155__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__A1 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A3 (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__A3 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A2 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A2 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__A4 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__B1 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A4 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A2 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__A2 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__I (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A1 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A1 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A1 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__A2 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__A2 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__A2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__A2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__A3 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A1 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5951__A1 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__A1 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A1 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A1 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A2 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A2 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__A2 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A1 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__A1 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A2 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A2 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__A3 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__I (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__A1 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8369__I (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8300__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__B1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__A2 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8250__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__A2 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A2 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__B (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A2 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A1 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__A1 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__A3 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__A2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__A2 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A2 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A2 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A2 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A2 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A2 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__A2 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__A1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__A1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__A1 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__B2 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__A2 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__B2 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__I (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__B2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__I (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A1 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__A1 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__A1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__A1 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8209__A1 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7237__A1 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__A1 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A1 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8210__A1 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7945__A3 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__B2 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__B2 (.I(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8014__A1 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__A1 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A1 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__A1 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A2 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__A2 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A3 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__A2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__A2 (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A2 (.I(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A2 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A2 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A1 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__A2 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A1 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__A1 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A1 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A1 (.I(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__B (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A1 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__I (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__B1 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__A3 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__I (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__A1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__A3 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8045__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8028__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__I (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__A1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__A2 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A2 (.I(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__A2 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__A2 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__A1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7370__A1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6267__I (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__A2 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__A2 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6142__A2 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__A1 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__A1 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__A3 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__A4 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__B1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A4 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__A2 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A2 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__B (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A3 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__A3 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__A3 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__A2 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__A2 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__B2 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8128__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__I (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__A1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__A1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__I (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__I (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__B (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A2 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__B (.I(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7465__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__I (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A2 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__A2 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6361__A1 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A1 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__B (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__A1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__A1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__B1 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A4 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__B (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6289__A1 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__A2 (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__A3 (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A2 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__A2 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__I (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__A1 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__A1 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__A1 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7671__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__A1 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A1 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__B (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__A2 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A2 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__A2 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A2 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6352__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A1 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__A1 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8357__A1 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__I (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A1 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A1 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__A2 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__A2 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A1 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__I (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__A1 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7408__A1 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__A1 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__A2 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__A1 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7474__A1 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A2 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__A2 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7673__B2 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__I (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A3 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__A3 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7467__A1 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__A1 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__A1 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__A1 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__A2 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A2 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__I (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__B (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__A1 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__A1 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__A1 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__A1 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__A2 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A1 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__A3 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8398__A1 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__A1 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__A1 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__I (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7580__A1 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6547__I (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__A1 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A1 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A2 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__A2 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__A2 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A2 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A2 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8449__A2 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8432__A2 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__A2 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A2 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7580__A3 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7552__A2 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__A3 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A2 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__A3 (.I(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__B (.I(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__A1 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8273__A1 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__A1 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__I (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8399__A1 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8358__A1 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__A1 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A3 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__A2 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8448__A1 (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7569__A1 (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__A1 (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__A1 (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__B1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__B1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__B1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__A2 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__I (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__B1 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7060__A3 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6690__I (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__I (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__I (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8014__B1 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__A2 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7709__A2 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__I (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__B1 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7657__A2 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6634__A2 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__I (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__A2 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__A2 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6631__A2 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__I (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__A2 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7612__A2 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7596__A2 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A2 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6871__A2 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__A2 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6596__I (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A3 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__I (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__I (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__A2 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__A2 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__I (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__A2 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer10_I (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7780__A3 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7619__I (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6575__I (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8036__A2 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__A2 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__A4 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__I (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7724__A2 (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7673__A2 (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__A2 (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__A2 (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__A2 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__A2 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__I (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__A3 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__A3 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__A3 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__A3 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__A2 (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__A2 (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__I (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A2 (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__A2 (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__I (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__A4 (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__A1 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__A1 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6658__A1 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__A1 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7716__A2 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__A2 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__A2 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6595__A2 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__B1 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7851__B1 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__A1 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__B2 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7851__B2 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__A2 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8038__A2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__A4 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7714__A3 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6600__A2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6666__A1 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6614__A1 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__A2 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__I (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__A2 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6604__A2 (.I(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__A2 (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__A2 (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__A2 (.I(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__A3 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__B1 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__B1 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__B1 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7708__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__I (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__B1 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__A2 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__A2 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__I (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__A2 (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__A2 (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__A2 (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__A2 (.I(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__C (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7822__A1 (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7115__I (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__A1 (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8016__A3 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7822__A3 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__A3 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__A2 (.I(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8107__A2 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7220__A2 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__A2 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6622__I (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8098__A2 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7645__A2 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__A2 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__I (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__A2 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__B1 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__I (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7658__A2 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7647__A2 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__A2 (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__I (.I(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__I (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6631__A4 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__A1 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__A1 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__A1 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6634__A1 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7945__B2 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__A2 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__A2 (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__I (.I(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7789__A2 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__A3 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7663__A2 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__I (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7581__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6638__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6689__A2 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6639__A2 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7029__A2 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__A2 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__A2 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__A2 (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__I (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6645__I (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__B1 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__A2 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__A4 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__A4 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7726__A2 (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__A2 (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6863__A2 (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__A2 (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__A2 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A2 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__A2 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__A2 (.I(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__A2 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__A4 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__A1 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__A2 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__A2 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7841__I (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A3 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__A3 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__A2 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__A2 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__A2 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__I (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6676__I (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8110__A2 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7208__A2 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__I (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__B1 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__A3 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7273__A2 (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__I (.I(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7696__A2 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__A2 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__A2 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6679__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7770__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7647__A3 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6682__A4 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6811__A1 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__A1 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__A1 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7929__A2 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7837__A2 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7059__A2 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__A2 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__A3 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__A3 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__A1 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__A1 (.I(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7591__A2 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__A2 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__A4 (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__I (.I(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__C (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__A3 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6747__A1 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__A1 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__B2 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6759__A1 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__A1 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7159__A1 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__A1 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__A1 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__A1 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__I (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__I (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7938__A2 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__A2 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__A2 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__A2 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__A3 (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__B1 (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__A3 (.I(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__B1 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__B1 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7719__B1 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6719__A1 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7717__A2 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6953__A2 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__A2 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__A2 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__B2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__B2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7719__B2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6719__A2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8134__A2 (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8045__A2 (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6720__A2 (.I(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__B1 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6759__A2 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__A2 (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6747__A2 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__A2 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__A3 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__A1 (.I(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7840__A2 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7107__A2 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__A2 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__I (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8111__A2 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7269__A2 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__I (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__I (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7991__A2 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7698__A2 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6791__A2 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__I (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__A2 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__A2 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6835__A2 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6754__A2 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__B2 (.I(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6782__A1 (.I(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8132__A2 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7793__A2 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__A2 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__A2 (.I(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6853__A1 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__B (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__A1 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__B2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8123__A2 (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__I (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6771__A2 (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7152__I (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__I (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6774__I (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7938__B1 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__A4 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__I (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__B1 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__A3 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__A1 (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__I (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8028__A4 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7028__A2 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__A2 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__A2 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6853__A3 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__A2 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6780__A2 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__B1 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6782__A2 (.I(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__A2 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__A2 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__A3 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6816__A2 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__A3 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6798__I (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__A1 (.I(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7108__A2 (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__A2 (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6801__I (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8089__A2 (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8010__A2 (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7270__A2 (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__I (.I(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8193__A2 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7924__A2 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A2 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6803__I (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8300__A2 (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8251__A2 (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__A2 (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6805__I (.I(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__A1 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6882__A1 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6898__A1 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__A1 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__A3 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6825__A1 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8250__A2 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7370__A2 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6999__I (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__A2 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6825__A2 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7824__A2 (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7346__A2 (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__A2 (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__A2 (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6899__A2 (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__A2 (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__A1 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6906__A1 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__A1 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6921__A1 (.I(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__A1 (.I(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7954__A2 (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7305__A2 (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__I (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__A2 (.I(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6921__A2 (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__A2 (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__A2 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__A2 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7020__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6855__I (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6846__I (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7789__B1 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__A4 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7663__B1 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__A2 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6917__A1 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__A1 (.I(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__A1 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__A1 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__A1 (.I(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8206__A2 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7667__A2 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__A3 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__I (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__A2 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__A2 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__A2 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__A1 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__A1 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7947__A2 (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7622__A2 (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__A3 (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__A3 (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7474__A2 (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__B1 (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__A4 (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__A1 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__A1 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__A1 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7028__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6863__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__A2 (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6862__I (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8276__A2 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8217__A2 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8044__A2 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6863__B1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__A2 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__A1 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__A2 (.I(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__B1 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__A2 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__A3 (.I(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__A2 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6946__A2 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__A2 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6871__B (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7060__A4 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7059__B1 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__I (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__I (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7721__A2 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__A2 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__A4 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__A2 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__A2 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__A2 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__A2 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__A3 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6917__A2 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__A2 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6895__A2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__A2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6882__A3 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6885__I (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__A1 (.I(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__A2 (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6888__I (.I(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8185__A2 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__A2 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__I (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__I (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7826__A2 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7425__A2 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__A2 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__I (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__I (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A1 (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__A1 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__A1 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__B2 (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__A1 (.I(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__A1 (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__A1 (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A2 (.I(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__A3 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6915__A2 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__A1 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__A1 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__A1 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__B2 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6936__A1 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8191__A2 (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8009__A2 (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7207__A2 (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__A2 (.I(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7052__A1 (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__A2 (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8013__A3 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__A3 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7063__A3 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__A3 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7061__A1 (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__A1 (.I(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__A1 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7273__B2 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__A1 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6933__A1 (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8274__A2 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7868__A2 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7127__I (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6933__A2 (.I(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__A3 (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7051__A2 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__A2 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__A3 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__A2 (.I(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6936__A2 (.I(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7010__A1 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__A1 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__A2 (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__A2 (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7013__A1 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__A1 (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__B (.I(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__I (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__A2 (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__A2 (.I(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__B2 (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__A1 (.I(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7025__A1 (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__A2 (.I(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__I (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6964__I (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8325__A2 (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__I (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__A4 (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__A2 (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7037__A2 (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7025__A2 (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__A3 (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7013__B (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__A3 (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__A3 (.I(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7010__A2 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__A2 (.I(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6992__A2 (.I(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6991__A2 (.I(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6971__A3 (.I(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__A2 (.I(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__A2 (.I(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A3 (.I(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__A2 (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6978__I (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__A1 (.I(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__I (.I(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__A2 (.I(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6979__I (.I(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8183__A2 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7277__A2 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__I (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8185__B1 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__B1 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__I (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6981__I (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8371__A2 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7987__A2 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7458__A1 (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6982__I (.I(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7077__A1 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__A1 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7759__A2 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__A2 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__A2 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__A2 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8255__A2 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7433__I (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__A2 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__A2 (.I(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7432__A2 (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A2 (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__I (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__A2 (.I(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7076__A2 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7008__A2 (.I(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7098__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__A1 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__A1 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7022__A1 (.I(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__A1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__A1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__A2 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__A3 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__B (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__A3 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__A2 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__A2 (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7031__A2 (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8216__A2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__A2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__B1 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__A2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7358__A3 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__A3 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__A3 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__A3 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__A1 (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__B (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__A2 (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__A2 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A3 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__A1 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7045__A1 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7418__I (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__I (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7358__A4 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__I (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__A2 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__A2 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7098__A2 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__A2 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__A2 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7087__A1 (.I(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__A1 (.I(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7102__A1 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__A1 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__A1 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__A1 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__A2 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7059__A1 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__A1 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7101__A1 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__A2 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__A1 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7111__A1 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__A2 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7957__A2 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__A4 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__I (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7065__A2 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7101__A2 (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7100__I (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__A3 (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7087__A2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__A2 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8302__A2 (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7994__A2 (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7909__A2 (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7084__A2 (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7178__A1 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7095__A1 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__A1 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__A3 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7183__A3 (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7093__A1 (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7177__A2 (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7094__A2 (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__A1 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__A1 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7184__A1 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__A1 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__B1 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__A2 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__A1 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A1 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__I (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A1 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__A1 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__I (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7121__A2 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8017__A1 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7838__A1 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7718__C (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__A1 (.I(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7928__A3 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__A3 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7710__A3 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__A3 (.I(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7184__A2 (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__A2 (.I(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A1 (.I(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__I (.I(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4419__I (.I(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__I (.I(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__A1 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__A1 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__A2 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8213__A2 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8046__A2 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__A2 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__A2 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7200__A1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7142__A1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7869__A2 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__A2 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7299__A2 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7136__A2 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7140__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A2 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A2 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__I (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__I (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__A1 (.I(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__I (.I(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8211__A2 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__A4 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7155__A2 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7153__A4 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7959__A2 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7290__A2 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7158__I (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7361__I (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7272__I (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7159__A2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__A2 (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__A2 (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__A3 (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A4 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__A4 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A3 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__A4 (.I(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7181__A2 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__A2 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__A3 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7253__A1 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7190__A1 (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__B2 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__A2 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__A2 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__A2 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__A1 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7245__A1 (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__A1 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7214__A1 (.I(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6871__A1 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__A1 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__I (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__A1 (.I(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7264__A1 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__A1 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7258__A2 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__A2 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__A1 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__B1 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__B1 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A1 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7262__A1 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7243__A1 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8030__A2 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7356__A2 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7304__A2 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7222__A2 (.I(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A2 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A1 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A2 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A1 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__A1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__A1 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7342__I (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__A1 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7232__A1 (.I(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7232__A2 (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__A1 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__A1 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7239__A1 (.I(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7354__A1 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__A1 (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__B (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__A2 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__A2 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7239__A2 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6606__A3 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__A2 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A3 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A2 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__A2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7316__A2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7247__A3 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__I (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A3 (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__I (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__I (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__I (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7389__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7329__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7328__A1 (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__A1 (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8172__A2 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7510__A2 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__A2 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__A2 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7330__A2 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__A2 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__A1 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__A1 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7333__A1 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7282__A1 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7434__A3 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7271__A2 (.I(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__A1 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7276__A1 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8031__A2 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__A2 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__A4 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7273__B1 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__A2 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7276__A2 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7394__A1 (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__A1 (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7280__A1 (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7280__A2 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7343__A2 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__A2 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__A1 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__A1 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7407__A1 (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7360__A1 (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7302__B (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7354__A2 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__A2 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__A1 (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__I (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__I (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7369__A1 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__A1 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7369__A2 (.I(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__A2 (.I(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__A1 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A1 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A1 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4298__I (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7387__A2 (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7382__A2 (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7319__A2 (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7388__A1 (.I(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7325__A1 (.I(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__A1 (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A1 (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__A1 (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A1 (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7388__A2 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7325__A2 (.I(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7394__A2 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__A2 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A1 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__I (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__A1 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__I (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7456__A1 (.I(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7426__A2 (.I(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__B (.I(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7427__A2 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7349__A2 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7401__A1 (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__A1 (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__A1 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__A1 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A1 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__A1 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7473__I (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7413__A1 (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7359__B (.I(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7407__A2 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7360__A2 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8280__A2 (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7514__I (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__I (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__A4 (.I(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7416__I (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7364__A1 (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7364__A2 (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__A2 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7366__A2 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__B2 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7374__A1 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__A1 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7373__A1 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__A1 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__A3 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__A4 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__A2 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7493__A1 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7442__A1 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7489__A1 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7440__A1 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7488__A1 (.I(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7439__A1 (.I(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A1 (.I(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7463__A1 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7414__A1 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7477__A4 (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7412__A1 (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__A3 (.I(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__A2 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__A2 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7479__I (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__A2 (.I(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7523__A1 (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7458__A2 (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7426__A3 (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7450__A1 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7437__A1 (.I(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__A2 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__A2 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__A2 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A1 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8303__A2 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7907__A2 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7465__A2 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7434__A2 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7449__A2 (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7436__A2 (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__I (.I(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__I (.I(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7532__A2 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7495__A2 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7446__A2 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__A1 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__A2 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__A1 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A2 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__C (.I(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7460__A1 (.I(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__A1 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7459__A1 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7523__A2 (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__A2 (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7459__A2 (.I(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7504__A1 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7484__A1 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8319__A2 (.I(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8181__A2 (.I(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8141__A2 (.I(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7467__A2 (.I(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__I (.I(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4314__I (.I(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__A1 (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7535__A1 (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7497__A2 (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__A3 (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__I (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__A2 (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__A1 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__A1 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__A1 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8400__A2 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8361__A2 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8352__I (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__A4 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__B (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__A2 (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__I (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__B (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__A1 (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__A1 (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__I (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7537__I (.I(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A1 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A1 (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4522__I (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__I (.I(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__B2 (.I(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A1 (.I(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A1 (.I(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A2 (.I(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7564__I (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7576__A1 (.I(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__A1 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__A1 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7615__A1 (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7595__A1 (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7582__A1 (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7582__A2 (.I(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A1 (.I(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A1 (.I(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__I (.I(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__I (.I(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__A1 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__A1 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__A2 (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__A2 (.I(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7594__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__A1 (.I(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__I (.I(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__A1 (.I(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__A1 (.I(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__A2 (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7594__A2 (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A1 (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__A1 (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__A2 (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__A2 (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7987__A1 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7909__A1 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7647__A1 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7610__I (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A3 (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__A3 (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__A3 (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__A3 (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__A2 (.I(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7865__A2 (.I(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7725__A2 (.I(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7620__A2 (.I(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__A1 (.I(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__A2 (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7663__B2 (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7622__A1 (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__A1 (.I(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__A2 (.I(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__A3 (.I(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7695__A2 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7656__A2 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__A2 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7626__A2 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7703__A2 (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7702__A2 (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7655__A2 (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7626__A3 (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A2 (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A2 (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4356__I (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__I (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A2 (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A2 (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A1 (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A1 (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7746__A1 (.I(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7734__A1 (.I(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__A1 (.I(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__A1 (.I(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__A1 (.I(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__A1 (.I(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__A1 (.I(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7753__A2 (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7697__A2 (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7660__A1 (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7695__A3 (.I(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7661__A2 (.I(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__A1 (.I(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7663__A1 (.I(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__A1 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__A2 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A1 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__I (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7706__A1 (.I(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7705__A1 (.I(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7675__A1 (.I(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7706__A2 (.I(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7705__A2 (.I(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7675__A2 (.I(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7724__A3 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7673__B1 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__A3 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7717__A1 (.I(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__B1 (.I(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__B1 (.I(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A2 (.I(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7703__A3 (.I(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7702__B (.I(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7676__A3 (.I(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A2 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A4 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A2 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A3 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7880__A1 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7743__A1 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7736__A1 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7742__A1 (.I(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7735__A1 (.I(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7745__A1 (.I(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7744__A1 (.I(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7734__A2 (.I(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7749__A1 (.I(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7701__A1 (.I(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7699__A2 (.I(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__I (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__I (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__I (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__I (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7766__A1 (.I(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__A1 (.I(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7731__A1 (.I(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7754__A2 (.I(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7712__A2 (.I(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7851__C (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__I (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__I (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__B (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7768__A1 (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7723__A1 (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__A1 (.I(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7852__B1 (.I(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7718__B1 (.I(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__A2 (.I(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7852__B2 (.I(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7718__B2 (.I(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7768__A2 (.I(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7723__A2 (.I(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__I (.I(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__I (.I(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7830__A1 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7777__A1 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__A1 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7728__A1 (.I(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7728__A2 (.I(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7776__A2 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7729__A2 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7750__A2 (.I(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__A2 (.I(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A1 (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__I (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__I (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__A1 (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__A1 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__B1 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__B1 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__A1 (.I(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7812__A1 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7803__A1 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A2 (.I(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__I (.I(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__A1 (.I(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7764__A1 (.I(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8014__A3 (.I(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7838__A3 (.I(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__A3 (.I(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__A3 (.I(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7819__A2 (.I(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7760__A2 (.I(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7813__A2 (.I(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__A2 (.I(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__B2 (.I(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__B2 (.I(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A2 (.I(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__A2 (.I(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7923__A1 (.I(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7833__A1 (.I(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__A1 (.I(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7905__A1 (.I(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7772__A2 (.I(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A2 (.I(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A2 (.I(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A2 (.I(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__B1 (.I(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7833__A2 (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__A2 (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7821__A2 (.I(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7775__A2 (.I(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7836__B2 (.I(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7786__A1 (.I(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7836__A1 (.I(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__A3 (.I(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__A1 (.I(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7864__A2 (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7835__A2 (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7834__A2 (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7785__A3 (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__A4 (.I(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7794__A1 (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7794__A2 (.I(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7847__I (.I(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7797__A2 (.I(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7934__A2 (.I(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7796__I (.I(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7831__B (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7799__A2 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7811__A2 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7802__A2 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__A1 (.I(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__I (.I(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__I (.I(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__A2 (.I(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__A1 (.I(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A1 (.I(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__A1 (.I(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7893__A1 (.I(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7877__A1 (.I(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__A1 (.I(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7829__A1 (.I(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7903__A1 (.I(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7843__A1 (.I(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7823__A2 (.I(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A2 (.I(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__A2 (.I(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__I (.I(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__A1 (.I(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7899__A1 (.I(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7825__A1 (.I(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7894__A2 (.I(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7828__A2 (.I(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A2 (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__I (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7902__A1 (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7846__A1 (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7901__A1 (.I(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7845__A1 (.I(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__A1 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7917__A1 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7844__A1 (.I(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8188__A3 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8017__A3 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7904__A3 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7842__A3 (.I(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7991__A3 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7903__A2 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7843__A3 (.I(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__A1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6908__A2 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__A1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__I (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7916__I (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7844__A2 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7901__A2 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7845__A2 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__A1 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7913__A1 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__A2 (.I(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7955__A1 (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7953__A1 (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7854__A1 (.I(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7955__A2 (.I(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7953__A2 (.I(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7854__A2 (.I(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7107__A1 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__I (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4352__I (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8040__I (.I(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__A1 (.I(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7861__A1 (.I(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7859__A2 (.I(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7947__A1 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__A1 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__B1 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7997__I (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__I (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7949__A1 (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7934__A3 (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7933__B1 (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7862__A1 (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A1 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__I (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A2 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__A1 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7872__A1 (.I(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__A1 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__B (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7920__A2 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7919__A2 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7872__A3 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7716__A1 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6595__A1 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__A1 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A1 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__A2 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7913__A2 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__A3 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7897__A2 (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7875__A2 (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7889__B2 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7878__A2 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A1 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__A1 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8067__A1 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7973__A1 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__A1 (.I(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__A1 (.I(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7982__A1 (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7912__A1 (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7981__A1 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7911__A1 (.I(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__A1 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7905__A2 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7981__A2 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7911__A2 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__A1 (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A2 (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__I (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A2 (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__A1 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__A1 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7921__A1 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8109__A1 (.I(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8096__A1 (.I(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7930__A1 (.I(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7923__A2 (.I(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__A2 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__A2 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7927__A1 (.I(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8090__A1 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__A2 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__A3 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7927__A2 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__B1 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7989__A2 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7932__A3 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7852__C (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7042__B (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__B (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__B (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8002__A1 (.I(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7963__A1 (.I(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__A2 (.I(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8028__A3 (.I(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__A3 (.I(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8029__A1 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7939__A2 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__A1 (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8022__A1 (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7998__A2 (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7949__A2 (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A1 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__I (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__B1 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8036__A3 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__A3 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8049__B (.I(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8035__A1 (.I(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7946__A1 (.I(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8035__A2 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7946__A2 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8035__A3 (.I(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__A3 (.I(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8007__A1 (.I(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7999__A1 (.I(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7962__A1 (.I(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__A2 (.I(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__I (.I(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A2 (.I(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4362__I (.I(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8006__A1 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7961__A1 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8141__A3 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8026__A2 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8025__A2 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__A2 (.I(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__A1 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__A1 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__I (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__A2 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__A2 (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__A2 (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__A2 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7967__A2 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A1 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A2 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__A2 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__A1 (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7996__A1 (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__A1 (.I(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8077__A1 (.I(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7996__A2 (.I(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__A2 (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8077__A2 (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7996__A3 (.I(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8088__B2 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8021__A1 (.I(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8088__A1 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__A1 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8021__A2 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8086__A1 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8085__A1 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8020__A1 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8108__A1 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8097__A2 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8018__A1 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8015__A2 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8189__A1 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8108__A2 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8018__A2 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8095__A1 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__A1 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__A1 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__B1 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__B1 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A1 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8094__A1 (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8093__A1 (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8059__A2 (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8102__A1 (.I(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8033__A1 (.I(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8182__A1 (.I(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8032__A1 (.I(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__A2 (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8041__A1 (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__A3 (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8041__A2 (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8128__A3 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8127__A1 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8053__S (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__A1 (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__A1 (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__I (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__I (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8055__A1 (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__I (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8062__A2 (.I(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A1 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A2 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A2 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A1 (.I(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A1 (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__A1 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8147__A1 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__A1 (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__A2 (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A1 (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__I (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8161__A1 (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8160__A1 (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8147__A2 (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8165__A1 (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8092__A1 (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__A1 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8091__A1 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__A2 (.I(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8091__A2 (.I(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8168__A1 (.I(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8146__A1 (.I(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__B1 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__A1 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__B1 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A2 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8167__A1 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8145__A1 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8171__A1 (.I(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8115__A1 (.I(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8170__A1 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8114__A1 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8106__A1 (.I(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8184__A1 (.I(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8172__B1 (.I(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__A2 (.I(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8180__A1 (.I(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8113__A1 (.I(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8112__A1 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8109__A2 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__I (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8113__A2 (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__A2 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__I (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__I (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8170__A2 (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8114__A2 (.I(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8175__A1 (.I(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8174__A1 (.I(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__A2 (.I(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__A1 (.I(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__A1 (.I(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8327__A2 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__A2 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8218__A2 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__A2 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A1 (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A1 (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__I (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__I (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8202__A1 (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8125__A1 (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__A1 (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__B (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8204__A1 (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8203__A1 (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8136__A2 (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8207__A1 (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8133__I0 (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__A2 (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__I (.I(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__A1 (.I(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A1 (.I(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__I (.I(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__A2 (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__A2 (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__A1 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A2 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__I (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A2 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8157__A3 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8156__B (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__A2 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8233__A1 (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8230__A1 (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8235__A1 (.I(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8228__A1 (.I(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8234__A1 (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8227__A1 (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8237__A2 (.I(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8173__A2 (.I(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6606__A1 (.I(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A1 (.I(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A1 (.I(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A1 (.I(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8241__A1 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__A1 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8240__A1 (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8197__A1 (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A3 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8292__A1 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8243__A1 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8186__A1 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8186__A2 (.I(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8192__A1 (.I(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8189__A2 (.I(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8247__A1 (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8195__A1 (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8301__A1 (.I(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8192__A2 (.I(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__A1 (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__B1 (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__I (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8247__A2 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8195__A2 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8240__A2 (.I(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8197__A2 (.I(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8262__A1 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8222__A1 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__A2 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__B1 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__B1 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A1 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__A1 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A1 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__A1 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__I (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8265__A2 (.I(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8215__A2 (.I(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__A1 (.I(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A1 (.I(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A1 (.I(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__I (.I(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7943__A1 (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A1 (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A1 (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__I (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8342__A1 (.I(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8290__A1 (.I(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8341__A1 (.I(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8289__A1 (.I(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7945__A1 (.I(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A1 (.I(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A1 (.I(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A1 (.I(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8297__A1 (.I(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8259__A1 (.I(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A2 (.I(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__A2 (.I(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__A3 (.I(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A3 (.I(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8372__A1 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8254__A2 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8297__A2 (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8259__A2 (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8295__A1 (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8294__A1 (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__A2 (.I(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__A1 (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A1 (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__A1 (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__I (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8313__A1 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8312__A1 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8283__A2 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8447__A2 (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8400__A1 (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8359__A1 (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8269__A1 (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8316__A1 (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8278__A1 (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__A2 (.I(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A2 (.I(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__A2 (.I(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A4 (.I(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8322__A2 (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8275__S (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8315__A2 (.I(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8281__A2 (.I(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__B1 (.I(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8293__I (.I(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__A1 (.I(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__I (.I(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__I (.I(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8345__A1 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8336__A1 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8379__B2 (.I(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8335__A1 (.I(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8379__A1 (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8334__A1 (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8304__A1 (.I(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8301__A2 (.I(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8368__A1 (.I(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8306__A1 (.I(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8372__B2 (.I(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8305__A1 (.I(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8424__A1 (.I(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8394__A1 (.I(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8391__A3 (.I(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8304__A2 (.I(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8310__A2 (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8309__A2 (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__A1 (.I(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__B2 (.I(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__A1 (.I(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__I (.I(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8348__A1 (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__A1 (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8396__A1 (.I(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8361__A1 (.I(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8355__A1 (.I(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8321__A1 (.I(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8356__A2 (.I(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8326__S (.I(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__A1 (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A1 (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A1 (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__I (.I(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__A2 (.I(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8340__A2 (.I(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8416__A2 (.I(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8385__A2 (.I(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8343__A2 (.I(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__A1 (.I(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A1 (.I(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__I (.I(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__A1 (.I(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A1 (.I(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8405__A1 (.I(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8364__A1 (.I(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8429__A1 (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__A1 (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8363__A1 (.I(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6953__A1 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__A2 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__B1 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__I (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8409__A2 (.I(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8367__A2 (.I(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer11_I (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__B1 (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A3 (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7781__C (.I(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__B (.I(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__B (.I(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__B (.I(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_rebuffer9_I (.I(_3604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A1 (.I(_3604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__A2 (.I(_3604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__I (.I(_3604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A2 (.I(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A1 (.I(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A1 (.I(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__I (.I(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A4 (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__B1 (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A1 (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__I (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8453__A1 (.I(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8452__A1 (.I(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8439__A1 (.I(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A1 (.I(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A2 (.I(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__I (.I(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__I (.I(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8553__A1 (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8442__I (.I(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__A1 (.I(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__I (.I(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8534__A2 (.I(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8504__A2 (.I(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__A2 (.I(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__A2 (.I(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8526__A2 (.I(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__S (.I(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8471__I (.I(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8470__I (.I(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__B1 (.I(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8490__A2 (.I(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__B1 (.I(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8477__A2 (.I(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8477__B (.I(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8506__I (.I(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__A2 (.I(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8484__A2 (.I(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8475__A2 (.I(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8550__B (.I(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8526__A1 (.I(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8482__I (.I(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8476__I (.I(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8540__A2 (.I(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8502__A2 (.I(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__C1 (.I(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8477__C (.I(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8538__S0 (.I(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8536__S0 (.I(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8498__A2 (.I(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__A1 (.I(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8509__S1 (.I(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__S1 (.I(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8498__A1 (.I(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__B (.I(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8552__A2 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8533__A2 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8511__A2 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8485__A2 (.I(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__A1 (.I(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A1 (.I(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8524__I (.I(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8522__S0 (.I(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8493__A1 (.I(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8484__A1 (.I(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__C1 (.I(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__B1 (.I(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8485__B1 (.I(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8551__B (.I(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8512__I (.I(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8503__C (.I(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8487__I (.I(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8553__A2 (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8520__A2 (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8491__A2 (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__A2 (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8492__A1 (.I(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8532__A1 (.I(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8517__A1 (.I(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8503__A1 (.I(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8494__I (.I(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8547__A1 (.I(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8542__A1 (.I(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8519__A2 (.I(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8497__A2 (.I(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__S (.I(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8541__S (.I(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8515__A2 (.I(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8497__B1 (.I(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8500__A1 (.I(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__B1 (.I(_3697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8503__B (.I(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A1 (.I(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__C (.I(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__C (.I(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__I (.I(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__A1 (.I(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8551__A1 (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8522__S1 (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8509__S0 (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__S0 (.I(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8510__I (.I(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8547__B (.I(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8542__B (.I(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8532__B (.I(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__A2 (.I(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__A2 (.I(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__I (.I(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A1 (.I(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A1 (.I(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8517__A3 (.I(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8548__A2 (.I(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8543__A2 (.I(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8529__S (.I(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8519__C (.I(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8521__A1 (.I(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8521__A2 (.I(_3716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8523__I (.I(_3717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__A1 (.I(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8545__A1 (.I(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8538__S1 (.I(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8536__S1 (.I(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8525__A1 (.I(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8530__I (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__A1 (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__I (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__A1 (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A2 (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8537__I (.I(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8539__I (.I(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__I (.I(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__I (.I(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8549__A1 (.I(_3737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8551__C (.I(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__B1 (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__B1 (.I(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__A1 (.I(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A2 (.I(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A2 (.I(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__A1 (.I(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A3 (.I(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__A3 (.I(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A3 (.I(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__I (.I(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__A2 (.I(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A3 (.I(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A2 (.I(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__A2 (.I(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__I (.I(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__I (.I(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__A1 (.I(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__I (.I(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A2 (.I(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A2 (.I(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__I (.I(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__I (.I(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__A2 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__A2 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A2 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__A2 (.I(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__B2 (.I(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__I (.I(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__I (.I(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__B2 (.I(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__B2 (.I(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__B2 (.I(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__B2 (.I(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__I (.I(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__I (.I(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A3 (.I(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__A1 (.I(_3758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__A1 (.I(_3758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__A1 (.I(_3758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__A1 (.I(_3758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__B (.I(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6586__A1 (.I(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__C (.I(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__I (.I(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__B (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__A2 (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__A1 (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__I (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A1 (.I(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__I (.I(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A2 (.I(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__I (.I(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A2 (.I(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A2 (.I(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__A2 (.I(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A2 (.I(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__B2 (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__B2 (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__B2 (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__B2 (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__I (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__I (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A2 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__I (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__A1 (.I(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__A1 (.I(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A3 (.I(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__A2 (.I(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A2 (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A2 (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__A2 (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A2 (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__B2 (.I(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__B2 (.I(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__B2 (.I(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__B2 (.I(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__I (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__I (.I(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__A1 (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A2 (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A1 (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__I (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__B2 (.I(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__A1 (.I(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__I (.I(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__A3 (.I(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__B2 (.I(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A1 (.I(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__A2 (.I(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__A2 (.I(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__A2 (.I(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__B (.I(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__I (.I(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__I (.I(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6908__A1 (.I(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__A2 (.I(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__A1 (.I(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__I (.I(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__A1 (.I(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A1 (.I(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A1 (.I(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__I (.I(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__I (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A1 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A2 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A1 (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__A2 (.I(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A2 (.I(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A2 (.I(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__I (.I(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A3 (.I(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A2 (.I(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A4 (.I(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A3 (.I(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__B2 (.I(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__B2 (.I(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__B2 (.I(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__I (.I(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__B2 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__B2 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__B2 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__B2 (.I(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7060__A1 (.I(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7059__B2 (.I(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__I (.I(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__A1 (.I(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6638__A1 (.I(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__A2 (.I(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A2 (.I(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__I (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__A2 (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A2 (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__A2 (.I(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__I (.I(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__B2 (.I(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__B2 (.I(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__B2 (.I(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__A2 (.I(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A2 (.I(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__I (.I(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__I (.I(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8462__A2 (.I(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__A2 (.I(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__A2 (.I(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A3 (.I(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7904__A1 (.I(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__A1 (.I(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6608__A1 (.I(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__I (.I(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7842__A1 (.I(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__A1 (.I(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__A1 (.I(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__I (.I(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__A1 (.I(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A1 (.I(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__B (.I(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A1 (.I(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8463__A2 (.I(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__A2 (.I(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__A3 (.I(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A2 (.I(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__A1 (.I(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__A1 (.I(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__B1 (.I(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__B1 (.I(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__A1 (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__I (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8459__A2 (.I(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A2 (.I(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A3 (.I(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A3 (.I(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A1 (.I(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__B2 (.I(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__A1 (.I(_3802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__B2 (.I(_3802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__B1 (.I(_3802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__A1 (.I(_3802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__I (.I(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A3 (.I(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__I (.I(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A1 (.I(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A1 (.I(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__A3 (.I(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__I (.I(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__A1 (.I(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__A1 (.I(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A3 (.I(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__A1 (.I(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__I (.I(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__I (.I(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__I (.I(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A1 (.I(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A2 (.I(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__A2 (.I(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__I (.I(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__I (.I(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__A1 (.I(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__I (.I(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A1 (.I(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__I (.I(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A1 (.I(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__A1 (.I(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A2 (.I(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__A1 (.I(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7290__A1 (.I(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7019__A1 (.I(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__I (.I(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7222__A1 (.I(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7136__A1 (.I(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A3 (.I(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__I (.I(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__A1 (.I(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__A2 (.I(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__I (.I(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__A2 (.I(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__A1 (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__A1 (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A1 (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__B1 (.I(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A1 (.I(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__I (.I(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A1 (.I(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7063__A1 (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__I (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__B (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__I (.I(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A1 (.I(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__A1 (.I(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__A1 (.I(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A2 (.I(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A2 (.I(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__I (.I(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__I (.I(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A2 (.I(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A2 (.I(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A2 (.I(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A3 (.I(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A1 (.I(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A2 (.I(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__A1 (.I(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__A3 (.I(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A2 (.I(_3826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__A1 (.I(_3826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4512__A1 (.I(_3826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__A2 (.I(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__A2 (.I(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__B2 (.I(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__B1 (.I(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__B1 (.I(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__I (.I(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__I (.I(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A1 (.I(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__I (.I(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A3 (.I(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__A1 (.I(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__A1 (.I(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6771__A1 (.I(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__I (.I(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__A2 (.I(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__A2 (.I(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__A3 (.I(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A1 (.I(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A1 (.I(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__A1 (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__I (.I(_3840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__I (.I(_3840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__I (.I(_3840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__A1 (.I(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A1 (.I(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A1 (.I(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A2 (.I(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__A1 (.I(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__I (.I(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A2 (.I(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A1 (.I(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__I (.I(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A1 (.I(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__I (.I(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A2 (.I(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A1 (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__A1 (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__A2 (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__A1 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__A2 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__I (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A1 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A1 (.I(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__A1 (.I(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A2 (.I(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__B2 (.I(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__A2 (.I(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7029__A1 (.I(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__I (.I(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__I (.I(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__A1 (.I(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__B (.I(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A3 (.I(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__A2 (.I(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A4 (.I(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__A3 (.I(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__I (.I(_3858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__I (.I(_3858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A2 (.I(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__B2 (.I(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__I (.I(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A1 (.I(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__A1 (.I(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__A2 (.I(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__A2 (.I(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__I (.I(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__A1 (.I(_3862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__A2 (.I(_3862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__I (.I(_3862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7207__A1 (.I(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A2 (.I(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A2 (.I(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__I (.I(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7270__A1 (.I(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6835__A1 (.I(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__I (.I(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A2 (.I(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__A1 (.I(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A1 (.I(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A2 (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__I (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__I (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A1 (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A1 (.I(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A1 (.I(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A2 (.I(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__A2 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A2 (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__I (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__I (.I(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A2 (.I(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__A1 (.I(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A2 (.I(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A1 (.I(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A2 (.I(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__A2 (.I(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__A1 (.I(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__I (.I(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__A2 (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7273__A1 (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A2 (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__I (.I(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7346__A1 (.I(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__I (.I(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A1 (.I(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__A2 (.I(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A1 (.I(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__A1 (.I(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__A1 (.I(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__I (.I(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__A1 (.I(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A1 (.I(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A1 (.I(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__B1 (.I(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__A1 (.I(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__A1 (.I(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__I (.I(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__B2 (.I(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4556__A2 (.I(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A3 (.I(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A2 (.I(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A2 (.I(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__A1 (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__I (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__A2 (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__A1 (.I(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7432__A1 (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__A1 (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A1 (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__I (.I(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__A1 (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6791__A1 (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__I (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__I (.I(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7084__A1 (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__A1 (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A2 (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A1 (.I(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__I (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__A1 (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__I (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A1 (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__A1 (.I(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__A1 (.I(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A2 (.I(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A1 (.I(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A2 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__B1 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__B1 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__I (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__A1 (.I(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__A1 (.I(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__B1 (.I(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A3 (.I(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__I (.I(_3896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__I (.I(_3896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__A2 (.I(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__A1 (.I(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A2 (.I(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__I (.I(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__B2 (.I(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A4 (.I(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A1 (.I(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__I (.I(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__A2 (.I(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__B2 (.I(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__I (.I(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__I (.I(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__A2 (.I(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__A1 (.I(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A2 (.I(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A2 (.I(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A1 (.I(_3902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__A1 (.I(_3902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__A1 (.I(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__I (.I(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__I (.I(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A1 (.I(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__A2 (.I(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A1 (.I(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__A2 (.I(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A2 (.I(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__A1 (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__I (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__I (.I(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7304__A1 (.I(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A1 (.I(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__I (.I(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A1 (.I(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A1 (.I(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__I (.I(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__I (.I(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__A1 (.I(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A1 (.I(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A3 (.I(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__I (.I(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A1 (.I(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__I (.I(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A2 (.I(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A2 (.I(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__A2 (.I(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A2 (.I(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8051__A1 (.I(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__A1 (.I(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__B2 (.I(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A2 (.I(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__I (.I(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__I (.I(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A3 (.I(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__I (.I(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A2 (.I(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__I (.I(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__A2 (.I(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7410__A2 (.I(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A2 (.I(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A4 (.I(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__I (.I(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__A1 (.I(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A1 (.I(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A1 (.I(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A1 (.I(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A1 (.I(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__I (.I(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__I (.I(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__I (.I(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A2 (.I(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A2 (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__A2 (.I(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__I (.I(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__A2 (.I(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__A2 (.I(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A3 (.I(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A2 (.I(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__A3 (.I(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__C (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A3 (.I(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A3 (.I(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A1 (.I(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__B (.I(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__B (.I(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__I (.I(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__I (.I(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8016__A1 (.I(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8013__A1 (.I(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__I (.I(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__I (.I(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A2 (.I(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A1 (.I(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__A1 (.I(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A1 (.I(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__A1 (.I(_3949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__I (.I(_3949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__I (.I(_3949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__A1 (.I(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A3 (.I(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A3 (.I(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A3 (.I(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__A1 (.I(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__I (.I(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A2 (.I(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A3 (.I(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__B1 (.I(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__I (.I(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A1 (.I(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A1 (.I(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A1 (.I(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__B2 (.I(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__I (.I(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__I (.I(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A2 (.I(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__A1 (.I(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__A1 (.I(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A3 (.I(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A3 (.I(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A2 (.I(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__B2 (.I(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__C (.I(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__A1 (.I(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__A1 (.I(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__I (.I(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__A1 (.I(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A1 (.I(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A1 (.I(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__A1 (.I(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__A1 (.I(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__A1 (.I(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__A1 (.I(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__A2 (.I(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A2 (.I(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__C (.I(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__A2 (.I(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__I (.I(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A3 (.I(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__I (.I(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__I (.I(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__A1 (.I(_3965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__A1 (.I(_3965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__I (.I(_3965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A1 (.I(_3965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6887__B2 (.I(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__B1 (.I(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__B1 (.I(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7291__A1 (.I(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__A1 (.I(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__I (.I(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7224__A1 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__A1 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__I (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A2 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__A1 (.I(_3970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A1 (.I(_3970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__A1 (.I(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6775__A1 (.I(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__A1 (.I(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__I (.I(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__A1 (.I(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__I (.I(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__A1 (.I(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__I (.I(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A1 (.I(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A1 (.I(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A1 (.I(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A1 (.I(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__B2 (.I(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__B2 (.I(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__B2 (.I(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A2 (.I(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__A1 (.I(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__A1 (.I(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__B2 (.I(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__I (.I(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A1 (.I(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__A1 (.I(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__B2 (.I(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__A1 (.I(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7020__A1 (.I(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__A3 (.I(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__I (.I(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__I (.I(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8460__A2 (.I(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A1 (.I(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__A2 (.I(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__A2 (.I(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7153__A1 (.I(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__A1 (.I(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A1 (.I(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__I (.I(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A1 (.I(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__A1 (.I(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A1 (.I(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__A1 (.I(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__A3 (.I(_3986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__A3 (.I(_3986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A2 (.I(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A2 (.I(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__B (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__B (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__B (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__I (.I(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__C (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__B (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A1 (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__I (.I(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8188__A1 (.I(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7928__A1 (.I(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__I (.I(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__I (.I(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__A1 (.I(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__A1 (.I(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A1 (.I(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__A1 (.I(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__A1 (.I(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__B2 (.I(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__A1 (.I(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A1 (.I(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7356__A1 (.I(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6961__A1 (.I(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__A2 (.I(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__I (.I(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__A1 (.I(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__A1 (.I(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__A2 (.I(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A3 (.I(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__A1 (.I(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__A1 (.I(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A1 (.I(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A1 (.I(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A1 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__A1 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__A2 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__B1 (.I(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__A1 (.I(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__A2 (.I(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A2 (.I(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__A2 (.I(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__A1 (.I(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__I (.I(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A2 (.I(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A2 (.I(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__A1 (.I(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__A1 (.I(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__I (.I(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A3 (.I(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6863__B2 (.I(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6720__A1 (.I(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A1 (.I(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__A1 (.I(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__I (.I(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__I (.I(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A2 (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__B2 (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A1 (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__A2 (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__B (.I(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__A3 (.I(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A3 (.I(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A1 (.I(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A1 (.I(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A1 (.I(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__A2 (.I(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A1 (.I(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A2 (.I(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__A1 (.I(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A2 (.I(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__A2 (.I(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__B2 (.I(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__I (.I(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__A1 (.I(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A1 (.I(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__A1 (.I(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A1 (.I(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__I (.I(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A1 (.I(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__A1 (.I(_4034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__I (.I(_4034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__I (.I(_4034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7510__A1 (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7220__A1 (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__A1 (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A2 (.I(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A3 (.I(_4036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__A2 (.I(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A2 (.I(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A1 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__B2 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A2 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A1 (.I(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__A1 (.I(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A1 (.I(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A2 (.I(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A2 (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__A2 (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A2 (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__A1 (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__A1 (.I(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A1 (.I(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__A1 (.I(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__I (.I(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__I (.I(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A3 (.I(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__A1 (.I(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A1 (.I(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__I (.I(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__A2 (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A2 (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__I (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A2 (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__B (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__A3 (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A3 (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7719__C (.I(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A1 (.I(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__I (.I(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A1 (.I(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A2 (.I(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__A2 (.I(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A2 (.I(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A2 (.I(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A3 (.I(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A1 (.I(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A2 (.I(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A2 (.I(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__A1 (.I(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__B2 (.I(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A1 (.I(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__A1 (.I(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__A1 (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A1 (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A1 (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__A2 (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__A1 (.I(_4071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__A1 (.I(_4071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__I (.I(_4071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__I (.I(_4071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__A1 (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A1 (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A1 (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__I (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__A1 (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A1 (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__B2 (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__A3 (.I(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__A1 (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__A1 (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6761__A1 (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A1 (.I(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__B2 (.I(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__B2 (.I(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__B2 (.I(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A2 (.I(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A2 (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A2 (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__A2 (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__B1 (.I(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A2 (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A2 (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__I (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__A2 (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__A2 (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A1 (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A2 (.I(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7305__A1 (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__I (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A4 (.I(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A1 (.I(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__A1 (.I(_4087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__I (.I(_4087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__B2 (.I(_4087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__I (.I(_4087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__B2 (.I(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__B2 (.I(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__B2 (.I(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__A1 (.I(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__A1 (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__I (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__I (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__I (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7358__A1 (.I(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7236__A1 (.I(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__A1 (.I(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__A1 (.I(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__A2 (.I(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__A2 (.I(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__I (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__I (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__I (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__I (.I(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A3 (.I(_4093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A3 (.I(_4093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__A3 (.I(_4093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__B1 (.I(_4093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A1 (.I(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A2 (.I(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__A3 (.I(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__A3 (.I(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A3 (.I(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A3 (.I(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__A2 (.I(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A2 (.I(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A3 (.I(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__A2 (.I(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__A2 (.I(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__I (.I(_4107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__A1 (.I(_4107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A1 (.I(_4107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__A2 (.I(_4107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7106__A1 (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__A1 (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__A1 (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__I (.I(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__A1 (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__A1 (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A1 (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__I (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__A1 (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6682__A1 (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6631__A1 (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__I (.I(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__A1 (.I(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A2 (.I(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__A3 (.I(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A2 (.I(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__A1 (.I(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__A1 (.I(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__A1 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A1 (.I(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5818__B2 (.I(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A2 (.I(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__A1 (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__A1 (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__A1 (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__A2 (.I(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7269__A1 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7208__A1 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6929__A1 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__A2 (.I(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__A1 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__A2 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__I (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A2 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__A1 (.I(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__A1 (.I(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__A2 (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__A2 (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__A2 (.I(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A2 (.I(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__A1 (.I(_4149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__A1 (.I(_4149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A2 (.I(_4149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__A1 (.I(_4150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__A2 (.I(_4150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__B1 (.I(_4150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A1 (.I(_4150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A1 (.I(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A2 (.I(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A3 (.I(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A1 (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A1 (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A1 (.I(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__A1 (.I(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__A1 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__A1 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6592__A1 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__A1 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__A1 (.I(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__A1 (.I(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__A1 (.I(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__A1 (.I(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A2 (.I(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__I (.I(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__A2 (.I(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A1 (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A1 (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A1 (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__A1 (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__A2 (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__A2 (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A2 (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__A2 (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A1 (.I(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__A1 (.I(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A1 (.I(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__A1 (.I(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A1 (.I(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__A1 (.I(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__A1 (.I(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A2 (.I(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__A1 (.I(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__I (.I(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__A1 (.I(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__B2 (.I(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__A1 (.I(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A3 (.I(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A2 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A1 (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__I (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A1 (.I(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__A1 (.I(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__A1 (.I(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__A2 (.I(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__A2 (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__A2 (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__A3 (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__A3 (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A3 (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__A3 (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A3 (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__A3 (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A3 (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A3 (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A4 (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__B1 (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A4 (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__I (.I(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__A3 (.I(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A3 (.I(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A3 (.I(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A1 (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A2 (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A2 (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__A2 (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A2 (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__A2 (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A2 (.I(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__A2 (.I(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A2 (.I(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__A2 (.I(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7202__A1 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__B2 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__A1 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__I (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__A1 (.I(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A2 (.I(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A1 (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A1 (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A1 (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__A2 (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__A1 (.I(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__A1 (.I(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__A1 (.I(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__C (.I(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A3 (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A1 (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__A1 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6754__A1 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__B2 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A2 (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A2 (.I(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__A2 (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A2 (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A2 (.I(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__A1 (.I(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__A1 (.I(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__I (.I(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__A2 (.I(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__B2 (.I(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A1 (.I(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A2 (.I(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__A1 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7065__A1 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__I (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__I (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__A1 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A1 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A2 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A3 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__B1 (.I(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A2 (.I(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A1 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A1 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A1 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A1 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A2 (.I(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A3 (.I(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__A2 (.I(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__A1 (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__A1 (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A1 (.I(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A1 (.I(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__A1 (.I(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A2 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__A2 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__A1 (.I(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A2 (.I(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A1 (.I(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__A1 (.I(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A1 (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__A1 (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__A2 (.I(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7727__A2 (.I(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__A3 (.I(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__A2 (.I(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__A2 (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__A2 (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__I (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A2 (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__A2 (.I(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A2 (.I(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__A2 (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A2 (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__B (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A1 (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__A1 (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__A1 (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__A2 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__A2 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__A1 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A1 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A1 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A1 (.I(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A2 (.I(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A2 (.I(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A2 (.I(_4273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A1 (.I(_4273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A2 (.I(_4273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A2 (.I(_4273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A3 (.I(_4274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A2 (.I(_4274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A1 (.I(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__B2 (.I(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A1 (.I(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A1 (.I(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__B (.I(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_Clock_I (.I(clknet_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_Clock_I (.I(clknet_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_Clock_I (.I(clknet_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_Clock_I (.I(clknet_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_Clock_I (.I(clknet_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_Clock_I (.I(clknet_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_Clock_I (.I(clknet_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_Clock_I (.I(clknet_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(reset));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__A1 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__A3 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A2 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__A2 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8468__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8465__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8473__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8464__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__A2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output16_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output23_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_1_0_Clock_I (.I(clknet_3_0_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_0_0_Clock_I (.I(clknet_3_0_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_3_0_Clock_I (.I(clknet_3_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_2_0_Clock_I (.I(clknet_3_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_5_0_Clock_I (.I(clknet_3_2_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_4_0_Clock_I (.I(clknet_3_2_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_7_0_Clock_I (.I(clknet_3_3_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_6_0_Clock_I (.I(clknet_3_3_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_9_0_Clock_I (.I(clknet_3_4_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_8_0_Clock_I (.I(clknet_3_4_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_11_0_Clock_I (.I(clknet_3_5_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_10_0_Clock_I (.I(clknet_3_5_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_13_0_Clock_I (.I(clknet_3_6_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_12_0_Clock_I (.I(clknet_3_6_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_15_0_Clock_I (.I(clknet_3_7_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_14_0_Clock_I (.I(clknet_3_7_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__CLK (.I(clknet_4_0_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__CLK (.I(clknet_4_0_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8566__CLK (.I(clknet_4_0_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8567__CLK (.I(clknet_4_0_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8595__CLK (.I(clknet_4_0_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8603__CLK (.I(clknet_4_0_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8605__CLK (.I(clknet_4_0_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8623__CLK (.I(clknet_4_0_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8624__CLK (.I(clknet_4_0_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8637__CLK (.I(clknet_4_0_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8640__CLK (.I(clknet_4_0_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8641__CLK (.I(clknet_4_0_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8642__CLK (.I(clknet_4_0_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8564__CLK (.I(clknet_4_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8575__CLK (.I(clknet_4_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__CLK (.I(clknet_4_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__CLK (.I(clknet_4_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__CLK (.I(clknet_4_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8587__CLK (.I(clknet_4_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8604__CLK (.I(clknet_4_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8606__CLK (.I(clknet_4_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8607__CLK (.I(clknet_4_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8611__CLK (.I(clknet_4_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8613__CLK (.I(clknet_4_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8615__CLK (.I(clknet_4_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8616__CLK (.I(clknet_4_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8619__CLK (.I(clknet_4_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8620__CLK (.I(clknet_4_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8621__CLK (.I(clknet_4_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8622__CLK (.I(clknet_4_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8636__CLK (.I(clknet_4_1_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8555__CLK (.I(clknet_4_2_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__CLK (.I(clknet_4_2_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8557__CLK (.I(clknet_4_2_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__CLK (.I(clknet_4_2_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8589__CLK (.I(clknet_4_2_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8590__CLK (.I(clknet_4_2_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8612__CLK (.I(clknet_4_2_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8625__CLK (.I(clknet_4_2_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8626__CLK (.I(clknet_4_2_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8639__CLK (.I(clknet_4_2_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8568__CLK (.I(clknet_4_3_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8569__CLK (.I(clknet_4_3_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8570__CLK (.I(clknet_4_3_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8572__CLK (.I(clknet_4_3_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8573__CLK (.I(clknet_4_3_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8574__CLK (.I(clknet_4_3_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8596__CLK (.I(clknet_4_3_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8597__CLK (.I(clknet_4_3_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8599__CLK (.I(clknet_4_3_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8601__CLK (.I(clknet_4_3_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8614__CLK (.I(clknet_4_3_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8581__CLK (.I(clknet_4_4_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8582__CLK (.I(clknet_4_4_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8583__CLK (.I(clknet_4_4_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__CLK (.I(clknet_4_4_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8653__CLK (.I(clknet_4_4_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8654__CLK (.I(clknet_4_4_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8670__CLK (.I(clknet_4_4_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8671__CLK (.I(clknet_4_4_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8672__CLK (.I(clknet_4_4_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8673__CLK (.I(clknet_4_4_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8674__CLK (.I(clknet_4_4_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8676__CLK (.I(clknet_4_4_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8675__CLK (.I(clknet_4_5_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8687__CLK (.I(clknet_4_5_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8688__CLK (.I(clknet_4_5_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8689__CLK (.I(clknet_4_5_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8690__CLK (.I(clknet_4_5_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8691__CLK (.I(clknet_4_5_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8692__CLK (.I(clknet_4_5_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8693__CLK (.I(clknet_4_5_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8571__CLK (.I(clknet_4_6_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8579__CLK (.I(clknet_4_6_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__CLK (.I(clknet_4_6_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8586__CLK (.I(clknet_4_6_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8656__CLK (.I(clknet_4_6_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8657__CLK (.I(clknet_4_6_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8658__CLK (.I(clknet_4_6_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8618__CLK (.I(clknet_4_7_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8659__CLK (.I(clknet_4_7_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8678__CLK (.I(clknet_4_7_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8679__CLK (.I(clknet_4_7_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8680__CLK (.I(clknet_4_7_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8681__CLK (.I(clknet_4_7_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8694__CLK (.I(clknet_4_7_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8695__CLK (.I(clknet_4_7_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8697__CLK (.I(clknet_4_7_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8558__CLK (.I(clknet_4_8_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__CLK (.I(clknet_4_8_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8627__CLK (.I(clknet_4_8_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8628__CLK (.I(clknet_4_8_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8629__CLK (.I(clknet_4_8_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8643__CLK (.I(clknet_4_8_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8644__CLK (.I(clknet_4_8_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8646__CLK (.I(clknet_4_8_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8591__CLK (.I(clknet_4_9_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8598__CLK (.I(clknet_4_9_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8600__CLK (.I(clknet_4_9_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8602__CLK (.I(clknet_4_9_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8617__CLK (.I(clknet_4_9_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8638__CLK (.I(clknet_4_9_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8645__CLK (.I(clknet_4_9_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8560__CLK (.I(clknet_4_10_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__CLK (.I(clknet_4_10_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8562__CLK (.I(clknet_4_10_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__CLK (.I(clknet_4_10_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8593__CLK (.I(clknet_4_10_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8594__CLK (.I(clknet_4_10_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8630__CLK (.I(clknet_4_10_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8631__CLK (.I(clknet_4_10_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8647__CLK (.I(clknet_4_10_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8608__CLK (.I(clknet_4_11_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8609__CLK (.I(clknet_4_11_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8610__CLK (.I(clknet_4_11_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8632__CLK (.I(clknet_4_11_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8633__CLK (.I(clknet_4_11_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8634__CLK (.I(clknet_4_11_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8635__CLK (.I(clknet_4_11_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8648__CLK (.I(clknet_4_11_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8649__CLK (.I(clknet_4_11_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8650__CLK (.I(clknet_4_11_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8651__CLK (.I(clknet_4_11_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8652__CLK (.I(clknet_4_11_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8682__CLK (.I(clknet_4_11_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8577__CLK (.I(clknet_4_12_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8655__CLK (.I(clknet_4_12_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8661__CLK (.I(clknet_4_12_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8677__CLK (.I(clknet_4_12_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8683__CLK (.I(clknet_4_12_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8684__CLK (.I(clknet_4_12_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8698__CLK (.I(clknet_4_12_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8685__CLK (.I(clknet_4_13_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8686__CLK (.I(clknet_4_13_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8696__CLK (.I(clknet_4_13_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8699__CLK (.I(clknet_4_13_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8700__CLK (.I(clknet_4_13_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8701__CLK (.I(clknet_4_13_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8702__CLK (.I(clknet_4_13_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8554__CLK (.I(clknet_4_14_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8660__CLK (.I(clknet_4_14_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8662__CLK (.I(clknet_4_14_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8663__CLK (.I(clknet_4_14_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8664__CLK (.I(clknet_4_15_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8665__CLK (.I(clknet_4_15_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8666__CLK (.I(clknet_4_15_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8667__CLK (.I(clknet_4_15_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8668__CLK (.I(clknet_4_15_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8669__CLK (.I(clknet_4_15_0_Clock));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7623__A2 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__A1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__B1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1577 ();
 assign done = net33;
endmodule

