VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO matrix_multiply
  CLASS BLOCK ;
  FOREIGN matrix_multiply ;
  ORIGIN 0.000 0.000 ;
  SIZE 700.000 BY 600.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 660.240 596.000 660.800 600.000 ;
    END
  END clk
  PIN execute
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 680.960 596.000 681.520 600.000 ;
    END
  END execute
  PIN input_val[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.080 596.000 80.640 600.000 ;
    END
  END input_val[0]
  PIN input_val[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 596.000 101.360 600.000 ;
    END
  END input_val[1]
  PIN input_val[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 121.520 596.000 122.080 600.000 ;
    END
  END input_val[2]
  PIN input_val[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 142.240 596.000 142.800 600.000 ;
    END
  END input_val[3]
  PIN input_val[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 162.960 596.000 163.520 600.000 ;
    END
  END input_val[4]
  PIN input_val[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 183.680 596.000 184.240 600.000 ;
    END
  END input_val[5]
  PIN input_val[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.400 596.000 204.960 600.000 ;
    END
  END input_val[6]
  PIN input_val[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 596.000 225.680 600.000 ;
    END
  END input_val[7]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 596.000 598.640 600.000 ;
    END
  END reset
  PIN result[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 245.840 596.000 246.400 600.000 ;
    END
  END result[0]
  PIN result[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 453.040 596.000 453.600 600.000 ;
    END
  END result[10]
  PIN result[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 473.760 596.000 474.320 600.000 ;
    END
  END result[11]
  PIN result[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 494.480 596.000 495.040 600.000 ;
    END
  END result[12]
  PIN result[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 515.200 596.000 515.760 600.000 ;
    END
  END result[13]
  PIN result[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 535.920 596.000 536.480 600.000 ;
    END
  END result[14]
  PIN result[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 556.640 596.000 557.200 600.000 ;
    END
  END result[15]
  PIN result[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 577.360 596.000 577.920 600.000 ;
    END
  END result[16]
  PIN result[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 266.560 596.000 267.120 600.000 ;
    END
  END result[1]
  PIN result[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 287.280 596.000 287.840 600.000 ;
    END
  END result[2]
  PIN result[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 308.000 596.000 308.560 600.000 ;
    END
  END result[3]
  PIN result[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 328.720 596.000 329.280 600.000 ;
    END
  END result[4]
  PIN result[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 349.440 596.000 350.000 600.000 ;
    END
  END result[5]
  PIN result[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 370.160 596.000 370.720 600.000 ;
    END
  END result[6]
  PIN result[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 390.880 596.000 391.440 600.000 ;
    END
  END result[7]
  PIN result[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 411.600 596.000 412.160 600.000 ;
    END
  END result[8]
  PIN result[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 432.320 596.000 432.880 600.000 ;
    END
  END result[9]
  PIN sel_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 17.920 596.000 18.480 600.000 ;
    END
  END sel_in[0]
  PIN sel_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 38.640 596.000 39.200 600.000 ;
    END
  END sel_in[1]
  PIN sel_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 596.000 59.920 600.000 ;
    END
  END sel_in[2]
  PIN sel_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 618.800 596.000 619.360 600.000 ;
    END
  END sel_out[0]
  PIN sel_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 639.520 596.000 640.080 600.000 ;
    END
  END sel_out[1]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 584.380 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 584.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 584.380 ;
    END
  END vssd1
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 693.280 585.050 ;
      LAYER Metal2 ;
        RECT 7.420 595.700 17.620 596.000 ;
        RECT 18.780 595.700 38.340 596.000 ;
        RECT 39.500 595.700 59.060 596.000 ;
        RECT 60.220 595.700 79.780 596.000 ;
        RECT 80.940 595.700 100.500 596.000 ;
        RECT 101.660 595.700 121.220 596.000 ;
        RECT 122.380 595.700 141.940 596.000 ;
        RECT 143.100 595.700 162.660 596.000 ;
        RECT 163.820 595.700 183.380 596.000 ;
        RECT 184.540 595.700 204.100 596.000 ;
        RECT 205.260 595.700 224.820 596.000 ;
        RECT 225.980 595.700 245.540 596.000 ;
        RECT 246.700 595.700 266.260 596.000 ;
        RECT 267.420 595.700 286.980 596.000 ;
        RECT 288.140 595.700 307.700 596.000 ;
        RECT 308.860 595.700 328.420 596.000 ;
        RECT 329.580 595.700 349.140 596.000 ;
        RECT 350.300 595.700 369.860 596.000 ;
        RECT 371.020 595.700 390.580 596.000 ;
        RECT 391.740 595.700 411.300 596.000 ;
        RECT 412.460 595.700 432.020 596.000 ;
        RECT 433.180 595.700 452.740 596.000 ;
        RECT 453.900 595.700 473.460 596.000 ;
        RECT 474.620 595.700 494.180 596.000 ;
        RECT 495.340 595.700 514.900 596.000 ;
        RECT 516.060 595.700 535.620 596.000 ;
        RECT 536.780 595.700 556.340 596.000 ;
        RECT 557.500 595.700 577.060 596.000 ;
        RECT 578.220 595.700 597.780 596.000 ;
        RECT 598.940 595.700 618.500 596.000 ;
        RECT 619.660 595.700 639.220 596.000 ;
        RECT 640.380 595.700 659.940 596.000 ;
        RECT 661.100 595.700 680.660 596.000 ;
        RECT 681.820 595.700 683.620 596.000 ;
        RECT 7.420 15.490 683.620 595.700 ;
      LAYER Metal3 ;
        RECT 7.370 15.540 682.550 587.860 ;
      LAYER Metal4 ;
        RECT 24.220 164.170 98.740 567.190 ;
        RECT 100.940 164.170 175.540 567.190 ;
        RECT 177.740 164.170 252.340 567.190 ;
        RECT 254.540 164.170 329.140 567.190 ;
        RECT 331.340 164.170 405.940 567.190 ;
        RECT 408.140 164.170 482.740 567.190 ;
        RECT 484.940 164.170 512.820 567.190 ;
  END
END matrix_multiply
END LIBRARY

