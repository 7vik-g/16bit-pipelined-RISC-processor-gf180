VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO io_interface
  CLASS BLOCK ;
  FOREIGN io_interface ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 1000.000 ;
  PIN clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 976.080 0.000 976.640 4.000 ;
    END
  END clk
  PIN data_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 638.960 996.000 639.520 1000.000 ;
    END
  END data_mem_addr[0]
  PIN data_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 649.040 996.000 649.600 1000.000 ;
    END
  END data_mem_addr[1]
  PIN data_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 659.120 996.000 659.680 1000.000 ;
    END
  END data_mem_addr[2]
  PIN data_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 669.200 996.000 669.760 1000.000 ;
    END
  END data_mem_addr[3]
  PIN data_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 679.280 996.000 679.840 1000.000 ;
    END
  END data_mem_addr[4]
  PIN data_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 689.360 996.000 689.920 1000.000 ;
    END
  END data_mem_addr[5]
  PIN data_mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 699.440 996.000 700.000 1000.000 ;
    END
  END data_mem_addr[6]
  PIN data_mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 709.520 996.000 710.080 1000.000 ;
    END
  END data_mem_addr[7]
  PIN data_read_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 642.320 996.000 642.880 1000.000 ;
    END
  END data_read_data[0]
  PIN data_read_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 733.040 996.000 733.600 1000.000 ;
    END
  END data_read_data[10]
  PIN data_read_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 739.760 996.000 740.320 1000.000 ;
    END
  END data_read_data[11]
  PIN data_read_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 746.480 996.000 747.040 1000.000 ;
    END
  END data_read_data[12]
  PIN data_read_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 753.200 996.000 753.760 1000.000 ;
    END
  END data_read_data[13]
  PIN data_read_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 759.920 996.000 760.480 1000.000 ;
    END
  END data_read_data[14]
  PIN data_read_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 766.640 996.000 767.200 1000.000 ;
    END
  END data_read_data[15]
  PIN data_read_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 652.400 996.000 652.960 1000.000 ;
    END
  END data_read_data[1]
  PIN data_read_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 662.480 996.000 663.040 1000.000 ;
    END
  END data_read_data[2]
  PIN data_read_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 672.560 996.000 673.120 1000.000 ;
    END
  END data_read_data[3]
  PIN data_read_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 682.640 996.000 683.200 1000.000 ;
    END
  END data_read_data[4]
  PIN data_read_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 692.720 996.000 693.280 1000.000 ;
    END
  END data_read_data[5]
  PIN data_read_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 702.800 996.000 703.360 1000.000 ;
    END
  END data_read_data[6]
  PIN data_read_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 712.880 996.000 713.440 1000.000 ;
    END
  END data_read_data[7]
  PIN data_read_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 719.600 996.000 720.160 1000.000 ;
    END
  END data_read_data[8]
  PIN data_read_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 726.320 996.000 726.880 1000.000 ;
    END
  END data_read_data[9]
  PIN data_write_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 645.680 996.000 646.240 1000.000 ;
    END
  END data_write_data[0]
  PIN data_write_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 736.400 996.000 736.960 1000.000 ;
    END
  END data_write_data[10]
  PIN data_write_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 743.120 996.000 743.680 1000.000 ;
    END
  END data_write_data[11]
  PIN data_write_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 749.840 996.000 750.400 1000.000 ;
    END
  END data_write_data[12]
  PIN data_write_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 756.560 996.000 757.120 1000.000 ;
    END
  END data_write_data[13]
  PIN data_write_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 763.280 996.000 763.840 1000.000 ;
    END
  END data_write_data[14]
  PIN data_write_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 770.000 996.000 770.560 1000.000 ;
    END
  END data_write_data[15]
  PIN data_write_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 655.760 996.000 656.320 1000.000 ;
    END
  END data_write_data[1]
  PIN data_write_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 665.840 996.000 666.400 1000.000 ;
    END
  END data_write_data[2]
  PIN data_write_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 675.920 996.000 676.480 1000.000 ;
    END
  END data_write_data[3]
  PIN data_write_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 686.000 996.000 686.560 1000.000 ;
    END
  END data_write_data[4]
  PIN data_write_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 696.080 996.000 696.640 1000.000 ;
    END
  END data_write_data[5]
  PIN data_write_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 706.160 996.000 706.720 1000.000 ;
    END
  END data_write_data[6]
  PIN data_write_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 716.240 996.000 716.800 1000.000 ;
    END
  END data_write_data[7]
  PIN data_write_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 722.960 996.000 723.520 1000.000 ;
    END
  END data_write_data[8]
  PIN data_write_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 729.680 996.000 730.240 1000.000 ;
    END
  END data_write_data[9]
  PIN dataw_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 635.600 996.000 636.160 1000.000 ;
    END
  END dataw_en
  PIN hlt
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 927.920 996.000 928.480 1000.000 ;
    END
  END hlt
  PIN instr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 776.720 996.000 777.280 1000.000 ;
    END
  END instr[0]
  PIN instr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 877.520 996.000 878.080 1000.000 ;
    END
  END instr[10]
  PIN instr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 887.600 996.000 888.160 1000.000 ;
    END
  END instr[11]
  PIN instr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 897.680 996.000 898.240 1000.000 ;
    END
  END instr[12]
  PIN instr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 907.760 996.000 908.320 1000.000 ;
    END
  END instr[13]
  PIN instr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 914.480 996.000 915.040 1000.000 ;
    END
  END instr[14]
  PIN instr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 921.200 996.000 921.760 1000.000 ;
    END
  END instr[15]
  PIN instr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 786.800 996.000 787.360 1000.000 ;
    END
  END instr[1]
  PIN instr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 796.880 996.000 797.440 1000.000 ;
    END
  END instr[2]
  PIN instr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 806.960 996.000 807.520 1000.000 ;
    END
  END instr[3]
  PIN instr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 817.040 996.000 817.600 1000.000 ;
    END
  END instr[4]
  PIN instr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 827.120 996.000 827.680 1000.000 ;
    END
  END instr[5]
  PIN instr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 837.200 996.000 837.760 1000.000 ;
    END
  END instr[6]
  PIN instr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 847.280 996.000 847.840 1000.000 ;
    END
  END instr[7]
  PIN instr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 857.360 996.000 857.920 1000.000 ;
    END
  END instr[8]
  PIN instr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 867.440 996.000 868.000 1000.000 ;
    END
  END instr[9]
  PIN instr_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 780.080 996.000 780.640 1000.000 ;
    END
  END instr_mem_addr[0]
  PIN instr_mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 880.880 996.000 881.440 1000.000 ;
    END
  END instr_mem_addr[10]
  PIN instr_mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 890.960 996.000 891.520 1000.000 ;
    END
  END instr_mem_addr[11]
  PIN instr_mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 901.040 996.000 901.600 1000.000 ;
    END
  END instr_mem_addr[12]
  PIN instr_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 790.160 996.000 790.720 1000.000 ;
    END
  END instr_mem_addr[1]
  PIN instr_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 800.240 996.000 800.800 1000.000 ;
    END
  END instr_mem_addr[2]
  PIN instr_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 810.320 996.000 810.880 1000.000 ;
    END
  END instr_mem_addr[3]
  PIN instr_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 820.400 996.000 820.960 1000.000 ;
    END
  END instr_mem_addr[4]
  PIN instr_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 830.480 996.000 831.040 1000.000 ;
    END
  END instr_mem_addr[5]
  PIN instr_mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 840.560 996.000 841.120 1000.000 ;
    END
  END instr_mem_addr[6]
  PIN instr_mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 850.640 996.000 851.200 1000.000 ;
    END
  END instr_mem_addr[7]
  PIN instr_mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 860.720 996.000 861.280 1000.000 ;
    END
  END instr_mem_addr[8]
  PIN instr_mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 870.800 996.000 871.360 1000.000 ;
    END
  END instr_mem_addr[9]
  PIN instr_write_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 783.440 996.000 784.000 1000.000 ;
    END
  END instr_write_data[0]
  PIN instr_write_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 884.240 996.000 884.800 1000.000 ;
    END
  END instr_write_data[10]
  PIN instr_write_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 894.320 996.000 894.880 1000.000 ;
    END
  END instr_write_data[11]
  PIN instr_write_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 904.400 996.000 904.960 1000.000 ;
    END
  END instr_write_data[12]
  PIN instr_write_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 911.120 996.000 911.680 1000.000 ;
    END
  END instr_write_data[13]
  PIN instr_write_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 917.840 996.000 918.400 1000.000 ;
    END
  END instr_write_data[14]
  PIN instr_write_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 924.560 996.000 925.120 1000.000 ;
    END
  END instr_write_data[15]
  PIN instr_write_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 793.520 996.000 794.080 1000.000 ;
    END
  END instr_write_data[1]
  PIN instr_write_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 803.600 996.000 804.160 1000.000 ;
    END
  END instr_write_data[2]
  PIN instr_write_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 813.680 996.000 814.240 1000.000 ;
    END
  END instr_write_data[3]
  PIN instr_write_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 823.760 996.000 824.320 1000.000 ;
    END
  END instr_write_data[4]
  PIN instr_write_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 833.840 996.000 834.400 1000.000 ;
    END
  END instr_write_data[5]
  PIN instr_write_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 843.920 996.000 844.480 1000.000 ;
    END
  END instr_write_data[6]
  PIN instr_write_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 854.000 996.000 854.560 1000.000 ;
    END
  END instr_write_data[7]
  PIN instr_write_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 864.080 996.000 864.640 1000.000 ;
    END
  END instr_write_data[8]
  PIN instr_write_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 874.160 996.000 874.720 1000.000 ;
    END
  END instr_write_data[9]
  PIN instrw_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 773.360 996.000 773.920 1000.000 ;
    END
  END instrw_en
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 71.120 996.000 71.680 1000.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.920 996.000 172.480 1000.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 182.000 996.000 182.560 1000.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 192.080 996.000 192.640 1000.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 202.160 996.000 202.720 1000.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 212.240 996.000 212.800 1000.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 222.320 996.000 222.880 1000.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 232.400 996.000 232.960 1000.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 242.480 996.000 243.040 1000.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 252.560 996.000 253.120 1000.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.640 996.000 263.200 1000.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 81.200 996.000 81.760 1000.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 272.720 996.000 273.280 1000.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 282.800 996.000 283.360 1000.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 292.880 996.000 293.440 1000.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 302.960 996.000 303.520 1000.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 313.040 996.000 313.600 1000.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 323.120 996.000 323.680 1000.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 333.200 996.000 333.760 1000.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 343.280 996.000 343.840 1000.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 353.360 996.000 353.920 1000.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 363.440 996.000 364.000 1000.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 91.280 996.000 91.840 1000.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 373.520 996.000 374.080 1000.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 383.600 996.000 384.160 1000.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 393.680 996.000 394.240 1000.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 403.760 996.000 404.320 1000.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 413.840 996.000 414.400 1000.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 423.920 996.000 424.480 1000.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 434.000 996.000 434.560 1000.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 444.080 996.000 444.640 1000.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 101.360 996.000 101.920 1000.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 111.440 996.000 112.000 1000.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 121.520 996.000 122.080 1000.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.600 996.000 132.160 1000.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 141.680 996.000 142.240 1000.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.760 996.000 152.320 1000.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.840 996.000 162.400 1000.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 74.480 996.000 75.040 1000.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 175.280 996.000 175.840 1000.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 185.360 996.000 185.920 1000.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 195.440 996.000 196.000 1000.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 205.520 996.000 206.080 1000.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.600 996.000 216.160 1000.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 225.680 996.000 226.240 1000.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 235.760 996.000 236.320 1000.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 245.840 996.000 246.400 1000.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.920 996.000 256.480 1000.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 266.000 996.000 266.560 1000.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.560 996.000 85.120 1000.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 276.080 996.000 276.640 1000.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 286.160 996.000 286.720 1000.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 296.240 996.000 296.800 1000.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 306.320 996.000 306.880 1000.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 316.400 996.000 316.960 1000.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 326.480 996.000 327.040 1000.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 336.560 996.000 337.120 1000.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 346.640 996.000 347.200 1000.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 356.720 996.000 357.280 1000.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 366.800 996.000 367.360 1000.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.640 996.000 95.200 1000.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 376.880 996.000 377.440 1000.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.960 996.000 387.520 1000.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 397.040 996.000 397.600 1000.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 407.120 996.000 407.680 1000.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 417.200 996.000 417.760 1000.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 427.280 996.000 427.840 1000.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 437.360 996.000 437.920 1000.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 447.440 996.000 448.000 1000.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.720 996.000 105.280 1000.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 114.800 996.000 115.360 1000.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.880 996.000 125.440 1000.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.960 996.000 135.520 1000.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 145.040 996.000 145.600 1000.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 155.120 996.000 155.680 1000.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 165.200 996.000 165.760 1000.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.840 996.000 78.400 1000.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 178.640 996.000 179.200 1000.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 188.720 996.000 189.280 1000.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 198.800 996.000 199.360 1000.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.880 996.000 209.440 1000.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.960 996.000 219.520 1000.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 229.040 996.000 229.600 1000.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 239.120 996.000 239.680 1000.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 249.200 996.000 249.760 1000.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 259.280 996.000 259.840 1000.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 269.360 996.000 269.920 1000.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.920 996.000 88.480 1000.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 279.440 996.000 280.000 1000.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 289.520 996.000 290.080 1000.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.600 996.000 300.160 1000.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 309.680 996.000 310.240 1000.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 319.760 996.000 320.320 1000.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.840 996.000 330.400 1000.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 339.920 996.000 340.480 1000.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 350.000 996.000 350.560 1000.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 360.080 996.000 360.640 1000.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 370.160 996.000 370.720 1000.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 98.000 996.000 98.560 1000.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 380.240 996.000 380.800 1000.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 390.320 996.000 390.880 1000.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 400.400 996.000 400.960 1000.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 410.480 996.000 411.040 1000.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 420.560 996.000 421.120 1000.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 430.640 996.000 431.200 1000.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 440.720 996.000 441.280 1000.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.800 996.000 451.360 1000.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 108.080 996.000 108.640 1000.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 118.160 996.000 118.720 1000.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 128.240 996.000 128.800 1000.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 138.320 996.000 138.880 1000.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 148.400 996.000 148.960 1000.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 158.480 996.000 159.040 1000.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.560 996.000 169.120 1000.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 954.240 0.000 954.800 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 961.520 0.000 962.080 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 968.800 0.000 969.360 4.000 ;
    END
  END irq[2]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.400 0.000 22.960 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 750.400 0.000 750.960 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 757.680 0.000 758.240 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 764.960 0.000 765.520 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 772.240 0.000 772.800 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 779.520 0.000 780.080 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 786.800 0.000 787.360 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 794.080 0.000 794.640 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 801.360 0.000 801.920 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 808.640 0.000 809.200 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 815.920 0.000 816.480 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 0.000 95.760 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 823.200 0.000 823.760 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 830.480 0.000 831.040 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 837.760 0.000 838.320 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 845.040 0.000 845.600 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 852.320 0.000 852.880 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 859.600 0.000 860.160 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 866.880 0.000 867.440 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 874.160 0.000 874.720 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 881.440 0.000 882.000 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 888.720 0.000 889.280 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 102.480 0.000 103.040 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 896.000 0.000 896.560 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 903.280 0.000 903.840 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 910.560 0.000 911.120 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 917.840 0.000 918.400 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 925.120 0.000 925.680 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 932.400 0.000 932.960 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 939.680 0.000 940.240 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 946.960 0.000 947.520 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 109.760 0.000 110.320 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.040 0.000 117.600 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.600 0.000 132.160 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 138.880 0.000 139.440 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 146.160 0.000 146.720 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 153.440 0.000 154.000 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 160.720 0.000 161.280 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.680 0.000 30.240 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 0.000 168.560 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 175.280 0.000 175.840 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 0.000 183.120 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 189.840 0.000 190.400 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 197.120 0.000 197.680 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.400 0.000 204.960 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 0.000 212.240 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 218.960 0.000 219.520 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 226.240 0.000 226.800 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 233.520 0.000 234.080 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 0.000 37.520 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 240.800 0.000 241.360 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.080 0.000 248.640 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 255.360 0.000 255.920 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.640 0.000 263.200 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 269.920 0.000 270.480 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 277.200 0.000 277.760 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 284.480 0.000 285.040 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 291.760 0.000 292.320 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 0.000 299.600 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 306.320 0.000 306.880 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 44.240 0.000 44.800 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 313.600 0.000 314.160 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 320.880 0.000 321.440 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 328.160 0.000 328.720 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 335.440 0.000 336.000 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 0.000 343.280 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 350.000 0.000 350.560 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 357.280 0.000 357.840 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 364.560 0.000 365.120 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 371.840 0.000 372.400 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 379.120 0.000 379.680 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 51.520 0.000 52.080 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 0.000 386.960 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 393.680 0.000 394.240 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 400.960 0.000 401.520 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 408.240 0.000 408.800 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 415.520 0.000 416.080 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 422.800 0.000 423.360 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 430.080 0.000 430.640 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 437.360 0.000 437.920 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 444.640 0.000 445.200 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 451.920 0.000 452.480 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 58.800 0.000 59.360 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 459.200 0.000 459.760 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 466.480 0.000 467.040 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 473.760 0.000 474.320 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 481.040 0.000 481.600 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 488.320 0.000 488.880 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 495.600 0.000 496.160 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 502.880 0.000 503.440 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 510.160 0.000 510.720 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 0.000 518.000 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 524.720 0.000 525.280 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 0.000 66.640 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 532.000 0.000 532.560 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 539.280 0.000 539.840 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 546.560 0.000 547.120 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 553.840 0.000 554.400 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 561.120 0.000 561.680 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 568.400 0.000 568.960 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 575.680 0.000 576.240 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 582.960 0.000 583.520 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 590.240 0.000 590.800 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 597.520 0.000 598.080 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.360 0.000 73.920 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 604.800 0.000 605.360 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 612.080 0.000 612.640 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 619.360 0.000 619.920 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 626.640 0.000 627.200 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 633.920 0.000 634.480 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 641.200 0.000 641.760 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 648.480 0.000 649.040 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 655.760 0.000 656.320 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 663.040 0.000 663.600 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 670.320 0.000 670.880 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 0.000 81.200 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 677.600 0.000 678.160 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 684.880 0.000 685.440 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 692.160 0.000 692.720 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 699.440 0.000 700.000 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 706.720 0.000 707.280 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 714.000 0.000 714.560 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 721.280 0.000 721.840 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 728.560 0.000 729.120 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 735.840 0.000 736.400 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 743.120 0.000 743.680 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.920 0.000 88.480 4.000 ;
    END
  END la_data_out[9]
  PIN reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 990.640 0.000 991.200 4.000 ;
    END
  END reset
  PIN start
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 983.360 0.000 983.920 4.000 ;
    END
  END start
  PIN uP_data_mem_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 457.520 996.000 458.080 1000.000 ;
    END
  END uP_data_mem_addr[0]
  PIN uP_data_mem_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 470.960 996.000 471.520 1000.000 ;
    END
  END uP_data_mem_addr[1]
  PIN uP_data_mem_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 484.400 996.000 484.960 1000.000 ;
    END
  END uP_data_mem_addr[2]
  PIN uP_data_mem_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 497.840 996.000 498.400 1000.000 ;
    END
  END uP_data_mem_addr[3]
  PIN uP_data_mem_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 511.280 996.000 511.840 1000.000 ;
    END
  END uP_data_mem_addr[4]
  PIN uP_data_mem_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 524.720 996.000 525.280 1000.000 ;
    END
  END uP_data_mem_addr[5]
  PIN uP_data_mem_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 538.160 996.000 538.720 1000.000 ;
    END
  END uP_data_mem_addr[6]
  PIN uP_data_mem_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 551.600 996.000 552.160 1000.000 ;
    END
  END uP_data_mem_addr[7]
  PIN uP_dataw_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 454.160 996.000 454.720 1000.000 ;
    END
  END uP_dataw_en
  PIN uP_instr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 460.880 996.000 461.440 1000.000 ;
    END
  END uP_instr[0]
  PIN uP_instr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 585.200 996.000 585.760 1000.000 ;
    END
  END uP_instr[10]
  PIN uP_instr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 595.280 996.000 595.840 1000.000 ;
    END
  END uP_instr[11]
  PIN uP_instr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 605.360 996.000 605.920 1000.000 ;
    END
  END uP_instr[12]
  PIN uP_instr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 615.440 996.000 616.000 1000.000 ;
    END
  END uP_instr[13]
  PIN uP_instr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 622.160 996.000 622.720 1000.000 ;
    END
  END uP_instr[14]
  PIN uP_instr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 628.880 996.000 629.440 1000.000 ;
    END
  END uP_instr[15]
  PIN uP_instr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 474.320 996.000 474.880 1000.000 ;
    END
  END uP_instr[1]
  PIN uP_instr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 487.760 996.000 488.320 1000.000 ;
    END
  END uP_instr[2]
  PIN uP_instr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 501.200 996.000 501.760 1000.000 ;
    END
  END uP_instr[3]
  PIN uP_instr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 514.640 996.000 515.200 1000.000 ;
    END
  END uP_instr[4]
  PIN uP_instr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 528.080 996.000 528.640 1000.000 ;
    END
  END uP_instr[5]
  PIN uP_instr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 541.520 996.000 542.080 1000.000 ;
    END
  END uP_instr[6]
  PIN uP_instr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 554.960 996.000 555.520 1000.000 ;
    END
  END uP_instr[7]
  PIN uP_instr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 565.040 996.000 565.600 1000.000 ;
    END
  END uP_instr[8]
  PIN uP_instr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 575.120 996.000 575.680 1000.000 ;
    END
  END uP_instr[9]
  PIN uP_instr_mem_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 464.240 996.000 464.800 1000.000 ;
    END
  END uP_instr_mem_addr[0]
  PIN uP_instr_mem_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 588.560 996.000 589.120 1000.000 ;
    END
  END uP_instr_mem_addr[10]
  PIN uP_instr_mem_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 598.640 996.000 599.200 1000.000 ;
    END
  END uP_instr_mem_addr[11]
  PIN uP_instr_mem_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 608.720 996.000 609.280 1000.000 ;
    END
  END uP_instr_mem_addr[12]
  PIN uP_instr_mem_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 477.680 996.000 478.240 1000.000 ;
    END
  END uP_instr_mem_addr[1]
  PIN uP_instr_mem_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 491.120 996.000 491.680 1000.000 ;
    END
  END uP_instr_mem_addr[2]
  PIN uP_instr_mem_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 504.560 996.000 505.120 1000.000 ;
    END
  END uP_instr_mem_addr[3]
  PIN uP_instr_mem_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 518.000 996.000 518.560 1000.000 ;
    END
  END uP_instr_mem_addr[4]
  PIN uP_instr_mem_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 531.440 996.000 532.000 1000.000 ;
    END
  END uP_instr_mem_addr[5]
  PIN uP_instr_mem_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 544.880 996.000 545.440 1000.000 ;
    END
  END uP_instr_mem_addr[6]
  PIN uP_instr_mem_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 558.320 996.000 558.880 1000.000 ;
    END
  END uP_instr_mem_addr[7]
  PIN uP_instr_mem_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 568.400 996.000 568.960 1000.000 ;
    END
  END uP_instr_mem_addr[8]
  PIN uP_instr_mem_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 578.480 996.000 579.040 1000.000 ;
    END
  END uP_instr_mem_addr[9]
  PIN uP_write_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 467.600 996.000 468.160 1000.000 ;
    END
  END uP_write_data[0]
  PIN uP_write_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 591.920 996.000 592.480 1000.000 ;
    END
  END uP_write_data[10]
  PIN uP_write_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 602.000 996.000 602.560 1000.000 ;
    END
  END uP_write_data[11]
  PIN uP_write_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 612.080 996.000 612.640 1000.000 ;
    END
  END uP_write_data[12]
  PIN uP_write_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 618.800 996.000 619.360 1000.000 ;
    END
  END uP_write_data[13]
  PIN uP_write_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 625.520 996.000 626.080 1000.000 ;
    END
  END uP_write_data[14]
  PIN uP_write_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 632.240 996.000 632.800 1000.000 ;
    END
  END uP_write_data[15]
  PIN uP_write_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 481.040 996.000 481.600 1000.000 ;
    END
  END uP_write_data[1]
  PIN uP_write_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 494.480 996.000 495.040 1000.000 ;
    END
  END uP_write_data[2]
  PIN uP_write_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 507.920 996.000 508.480 1000.000 ;
    END
  END uP_write_data[3]
  PIN uP_write_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 521.360 996.000 521.920 1000.000 ;
    END
  END uP_write_data[4]
  PIN uP_write_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 534.800 996.000 535.360 1000.000 ;
    END
  END uP_write_data[5]
  PIN uP_write_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 548.240 996.000 548.800 1000.000 ;
    END
  END uP_write_data[6]
  PIN uP_write_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 561.680 996.000 562.240 1000.000 ;
    END
  END uP_write_data[7]
  PIN uP_write_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 571.760 996.000 572.320 1000.000 ;
    END
  END uP_write_data[8]
  PIN uP_write_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 581.840 996.000 582.400 1000.000 ;
    END
  END uP_write_data[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 984.220 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 984.220 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 7.840 0.000 8.400 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 15.120 0.000 15.680 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 8.550 992.880 984.220 ;
      LAYER Metal2 ;
        RECT 7.980 995.700 70.820 999.510 ;
        RECT 71.980 995.700 74.180 999.510 ;
        RECT 75.340 995.700 77.540 999.510 ;
        RECT 78.700 995.700 80.900 999.510 ;
        RECT 82.060 995.700 84.260 999.510 ;
        RECT 85.420 995.700 87.620 999.510 ;
        RECT 88.780 995.700 90.980 999.510 ;
        RECT 92.140 995.700 94.340 999.510 ;
        RECT 95.500 995.700 97.700 999.510 ;
        RECT 98.860 995.700 101.060 999.510 ;
        RECT 102.220 995.700 104.420 999.510 ;
        RECT 105.580 995.700 107.780 999.510 ;
        RECT 108.940 995.700 111.140 999.510 ;
        RECT 112.300 995.700 114.500 999.510 ;
        RECT 115.660 995.700 117.860 999.510 ;
        RECT 119.020 995.700 121.220 999.510 ;
        RECT 122.380 995.700 124.580 999.510 ;
        RECT 125.740 995.700 127.940 999.510 ;
        RECT 129.100 995.700 131.300 999.510 ;
        RECT 132.460 995.700 134.660 999.510 ;
        RECT 135.820 995.700 138.020 999.510 ;
        RECT 139.180 995.700 141.380 999.510 ;
        RECT 142.540 995.700 144.740 999.510 ;
        RECT 145.900 995.700 148.100 999.510 ;
        RECT 149.260 995.700 151.460 999.510 ;
        RECT 152.620 995.700 154.820 999.510 ;
        RECT 155.980 995.700 158.180 999.510 ;
        RECT 159.340 995.700 161.540 999.510 ;
        RECT 162.700 995.700 164.900 999.510 ;
        RECT 166.060 995.700 168.260 999.510 ;
        RECT 169.420 995.700 171.620 999.510 ;
        RECT 172.780 995.700 174.980 999.510 ;
        RECT 176.140 995.700 178.340 999.510 ;
        RECT 179.500 995.700 181.700 999.510 ;
        RECT 182.860 995.700 185.060 999.510 ;
        RECT 186.220 995.700 188.420 999.510 ;
        RECT 189.580 995.700 191.780 999.510 ;
        RECT 192.940 995.700 195.140 999.510 ;
        RECT 196.300 995.700 198.500 999.510 ;
        RECT 199.660 995.700 201.860 999.510 ;
        RECT 203.020 995.700 205.220 999.510 ;
        RECT 206.380 995.700 208.580 999.510 ;
        RECT 209.740 995.700 211.940 999.510 ;
        RECT 213.100 995.700 215.300 999.510 ;
        RECT 216.460 995.700 218.660 999.510 ;
        RECT 219.820 995.700 222.020 999.510 ;
        RECT 223.180 995.700 225.380 999.510 ;
        RECT 226.540 995.700 228.740 999.510 ;
        RECT 229.900 995.700 232.100 999.510 ;
        RECT 233.260 995.700 235.460 999.510 ;
        RECT 236.620 995.700 238.820 999.510 ;
        RECT 239.980 995.700 242.180 999.510 ;
        RECT 243.340 995.700 245.540 999.510 ;
        RECT 246.700 995.700 248.900 999.510 ;
        RECT 250.060 995.700 252.260 999.510 ;
        RECT 253.420 995.700 255.620 999.510 ;
        RECT 256.780 995.700 258.980 999.510 ;
        RECT 260.140 995.700 262.340 999.510 ;
        RECT 263.500 995.700 265.700 999.510 ;
        RECT 266.860 995.700 269.060 999.510 ;
        RECT 270.220 995.700 272.420 999.510 ;
        RECT 273.580 995.700 275.780 999.510 ;
        RECT 276.940 995.700 279.140 999.510 ;
        RECT 280.300 995.700 282.500 999.510 ;
        RECT 283.660 995.700 285.860 999.510 ;
        RECT 287.020 995.700 289.220 999.510 ;
        RECT 290.380 995.700 292.580 999.510 ;
        RECT 293.740 995.700 295.940 999.510 ;
        RECT 297.100 995.700 299.300 999.510 ;
        RECT 300.460 995.700 302.660 999.510 ;
        RECT 303.820 995.700 306.020 999.510 ;
        RECT 307.180 995.700 309.380 999.510 ;
        RECT 310.540 995.700 312.740 999.510 ;
        RECT 313.900 995.700 316.100 999.510 ;
        RECT 317.260 995.700 319.460 999.510 ;
        RECT 320.620 995.700 322.820 999.510 ;
        RECT 323.980 995.700 326.180 999.510 ;
        RECT 327.340 995.700 329.540 999.510 ;
        RECT 330.700 995.700 332.900 999.510 ;
        RECT 334.060 995.700 336.260 999.510 ;
        RECT 337.420 995.700 339.620 999.510 ;
        RECT 340.780 995.700 342.980 999.510 ;
        RECT 344.140 995.700 346.340 999.510 ;
        RECT 347.500 995.700 349.700 999.510 ;
        RECT 350.860 995.700 353.060 999.510 ;
        RECT 354.220 995.700 356.420 999.510 ;
        RECT 357.580 995.700 359.780 999.510 ;
        RECT 360.940 995.700 363.140 999.510 ;
        RECT 364.300 995.700 366.500 999.510 ;
        RECT 367.660 995.700 369.860 999.510 ;
        RECT 371.020 995.700 373.220 999.510 ;
        RECT 374.380 995.700 376.580 999.510 ;
        RECT 377.740 995.700 379.940 999.510 ;
        RECT 381.100 995.700 383.300 999.510 ;
        RECT 384.460 995.700 386.660 999.510 ;
        RECT 387.820 995.700 390.020 999.510 ;
        RECT 391.180 995.700 393.380 999.510 ;
        RECT 394.540 995.700 396.740 999.510 ;
        RECT 397.900 995.700 400.100 999.510 ;
        RECT 401.260 995.700 403.460 999.510 ;
        RECT 404.620 995.700 406.820 999.510 ;
        RECT 407.980 995.700 410.180 999.510 ;
        RECT 411.340 995.700 413.540 999.510 ;
        RECT 414.700 995.700 416.900 999.510 ;
        RECT 418.060 995.700 420.260 999.510 ;
        RECT 421.420 995.700 423.620 999.510 ;
        RECT 424.780 995.700 426.980 999.510 ;
        RECT 428.140 995.700 430.340 999.510 ;
        RECT 431.500 995.700 433.700 999.510 ;
        RECT 434.860 995.700 437.060 999.510 ;
        RECT 438.220 995.700 440.420 999.510 ;
        RECT 441.580 995.700 443.780 999.510 ;
        RECT 444.940 995.700 447.140 999.510 ;
        RECT 448.300 995.700 450.500 999.510 ;
        RECT 451.660 995.700 453.860 999.510 ;
        RECT 455.020 995.700 457.220 999.510 ;
        RECT 458.380 995.700 460.580 999.510 ;
        RECT 461.740 995.700 463.940 999.510 ;
        RECT 465.100 995.700 467.300 999.510 ;
        RECT 468.460 995.700 470.660 999.510 ;
        RECT 471.820 995.700 474.020 999.510 ;
        RECT 475.180 995.700 477.380 999.510 ;
        RECT 478.540 995.700 480.740 999.510 ;
        RECT 481.900 995.700 484.100 999.510 ;
        RECT 485.260 995.700 487.460 999.510 ;
        RECT 488.620 995.700 490.820 999.510 ;
        RECT 491.980 995.700 494.180 999.510 ;
        RECT 495.340 995.700 497.540 999.510 ;
        RECT 498.700 995.700 500.900 999.510 ;
        RECT 502.060 995.700 504.260 999.510 ;
        RECT 505.420 995.700 507.620 999.510 ;
        RECT 508.780 995.700 510.980 999.510 ;
        RECT 512.140 995.700 514.340 999.510 ;
        RECT 515.500 995.700 517.700 999.510 ;
        RECT 518.860 995.700 521.060 999.510 ;
        RECT 522.220 995.700 524.420 999.510 ;
        RECT 525.580 995.700 527.780 999.510 ;
        RECT 528.940 995.700 531.140 999.510 ;
        RECT 532.300 995.700 534.500 999.510 ;
        RECT 535.660 995.700 537.860 999.510 ;
        RECT 539.020 995.700 541.220 999.510 ;
        RECT 542.380 995.700 544.580 999.510 ;
        RECT 545.740 995.700 547.940 999.510 ;
        RECT 549.100 995.700 551.300 999.510 ;
        RECT 552.460 995.700 554.660 999.510 ;
        RECT 555.820 995.700 558.020 999.510 ;
        RECT 559.180 995.700 561.380 999.510 ;
        RECT 562.540 995.700 564.740 999.510 ;
        RECT 565.900 995.700 568.100 999.510 ;
        RECT 569.260 995.700 571.460 999.510 ;
        RECT 572.620 995.700 574.820 999.510 ;
        RECT 575.980 995.700 578.180 999.510 ;
        RECT 579.340 995.700 581.540 999.510 ;
        RECT 582.700 995.700 584.900 999.510 ;
        RECT 586.060 995.700 588.260 999.510 ;
        RECT 589.420 995.700 591.620 999.510 ;
        RECT 592.780 995.700 594.980 999.510 ;
        RECT 596.140 995.700 598.340 999.510 ;
        RECT 599.500 995.700 601.700 999.510 ;
        RECT 602.860 995.700 605.060 999.510 ;
        RECT 606.220 995.700 608.420 999.510 ;
        RECT 609.580 995.700 611.780 999.510 ;
        RECT 612.940 995.700 615.140 999.510 ;
        RECT 616.300 995.700 618.500 999.510 ;
        RECT 619.660 995.700 621.860 999.510 ;
        RECT 623.020 995.700 625.220 999.510 ;
        RECT 626.380 995.700 628.580 999.510 ;
        RECT 629.740 995.700 631.940 999.510 ;
        RECT 633.100 995.700 635.300 999.510 ;
        RECT 636.460 995.700 638.660 999.510 ;
        RECT 639.820 995.700 642.020 999.510 ;
        RECT 643.180 995.700 645.380 999.510 ;
        RECT 646.540 995.700 648.740 999.510 ;
        RECT 649.900 995.700 652.100 999.510 ;
        RECT 653.260 995.700 655.460 999.510 ;
        RECT 656.620 995.700 658.820 999.510 ;
        RECT 659.980 995.700 662.180 999.510 ;
        RECT 663.340 995.700 665.540 999.510 ;
        RECT 666.700 995.700 668.900 999.510 ;
        RECT 670.060 995.700 672.260 999.510 ;
        RECT 673.420 995.700 675.620 999.510 ;
        RECT 676.780 995.700 678.980 999.510 ;
        RECT 680.140 995.700 682.340 999.510 ;
        RECT 683.500 995.700 685.700 999.510 ;
        RECT 686.860 995.700 689.060 999.510 ;
        RECT 690.220 995.700 692.420 999.510 ;
        RECT 693.580 995.700 695.780 999.510 ;
        RECT 696.940 995.700 699.140 999.510 ;
        RECT 700.300 995.700 702.500 999.510 ;
        RECT 703.660 995.700 705.860 999.510 ;
        RECT 707.020 995.700 709.220 999.510 ;
        RECT 710.380 995.700 712.580 999.510 ;
        RECT 713.740 995.700 715.940 999.510 ;
        RECT 717.100 995.700 719.300 999.510 ;
        RECT 720.460 995.700 722.660 999.510 ;
        RECT 723.820 995.700 726.020 999.510 ;
        RECT 727.180 995.700 729.380 999.510 ;
        RECT 730.540 995.700 732.740 999.510 ;
        RECT 733.900 995.700 736.100 999.510 ;
        RECT 737.260 995.700 739.460 999.510 ;
        RECT 740.620 995.700 742.820 999.510 ;
        RECT 743.980 995.700 746.180 999.510 ;
        RECT 747.340 995.700 749.540 999.510 ;
        RECT 750.700 995.700 752.900 999.510 ;
        RECT 754.060 995.700 756.260 999.510 ;
        RECT 757.420 995.700 759.620 999.510 ;
        RECT 760.780 995.700 762.980 999.510 ;
        RECT 764.140 995.700 766.340 999.510 ;
        RECT 767.500 995.700 769.700 999.510 ;
        RECT 770.860 995.700 773.060 999.510 ;
        RECT 774.220 995.700 776.420 999.510 ;
        RECT 777.580 995.700 779.780 999.510 ;
        RECT 780.940 995.700 783.140 999.510 ;
        RECT 784.300 995.700 786.500 999.510 ;
        RECT 787.660 995.700 789.860 999.510 ;
        RECT 791.020 995.700 793.220 999.510 ;
        RECT 794.380 995.700 796.580 999.510 ;
        RECT 797.740 995.700 799.940 999.510 ;
        RECT 801.100 995.700 803.300 999.510 ;
        RECT 804.460 995.700 806.660 999.510 ;
        RECT 807.820 995.700 810.020 999.510 ;
        RECT 811.180 995.700 813.380 999.510 ;
        RECT 814.540 995.700 816.740 999.510 ;
        RECT 817.900 995.700 820.100 999.510 ;
        RECT 821.260 995.700 823.460 999.510 ;
        RECT 824.620 995.700 826.820 999.510 ;
        RECT 827.980 995.700 830.180 999.510 ;
        RECT 831.340 995.700 833.540 999.510 ;
        RECT 834.700 995.700 836.900 999.510 ;
        RECT 838.060 995.700 840.260 999.510 ;
        RECT 841.420 995.700 843.620 999.510 ;
        RECT 844.780 995.700 846.980 999.510 ;
        RECT 848.140 995.700 850.340 999.510 ;
        RECT 851.500 995.700 853.700 999.510 ;
        RECT 854.860 995.700 857.060 999.510 ;
        RECT 858.220 995.700 860.420 999.510 ;
        RECT 861.580 995.700 863.780 999.510 ;
        RECT 864.940 995.700 867.140 999.510 ;
        RECT 868.300 995.700 870.500 999.510 ;
        RECT 871.660 995.700 873.860 999.510 ;
        RECT 875.020 995.700 877.220 999.510 ;
        RECT 878.380 995.700 880.580 999.510 ;
        RECT 881.740 995.700 883.940 999.510 ;
        RECT 885.100 995.700 887.300 999.510 ;
        RECT 888.460 995.700 890.660 999.510 ;
        RECT 891.820 995.700 894.020 999.510 ;
        RECT 895.180 995.700 897.380 999.510 ;
        RECT 898.540 995.700 900.740 999.510 ;
        RECT 901.900 995.700 904.100 999.510 ;
        RECT 905.260 995.700 907.460 999.510 ;
        RECT 908.620 995.700 910.820 999.510 ;
        RECT 911.980 995.700 914.180 999.510 ;
        RECT 915.340 995.700 917.540 999.510 ;
        RECT 918.700 995.700 920.900 999.510 ;
        RECT 922.060 995.700 924.260 999.510 ;
        RECT 925.420 995.700 927.620 999.510 ;
        RECT 928.780 995.700 991.620 999.510 ;
        RECT 7.980 4.300 991.620 995.700 ;
        RECT 8.700 3.500 14.820 4.300 ;
        RECT 15.980 3.500 22.100 4.300 ;
        RECT 23.260 3.500 29.380 4.300 ;
        RECT 30.540 3.500 36.660 4.300 ;
        RECT 37.820 3.500 43.940 4.300 ;
        RECT 45.100 3.500 51.220 4.300 ;
        RECT 52.380 3.500 58.500 4.300 ;
        RECT 59.660 3.500 65.780 4.300 ;
        RECT 66.940 3.500 73.060 4.300 ;
        RECT 74.220 3.500 80.340 4.300 ;
        RECT 81.500 3.500 87.620 4.300 ;
        RECT 88.780 3.500 94.900 4.300 ;
        RECT 96.060 3.500 102.180 4.300 ;
        RECT 103.340 3.500 109.460 4.300 ;
        RECT 110.620 3.500 116.740 4.300 ;
        RECT 117.900 3.500 124.020 4.300 ;
        RECT 125.180 3.500 131.300 4.300 ;
        RECT 132.460 3.500 138.580 4.300 ;
        RECT 139.740 3.500 145.860 4.300 ;
        RECT 147.020 3.500 153.140 4.300 ;
        RECT 154.300 3.500 160.420 4.300 ;
        RECT 161.580 3.500 167.700 4.300 ;
        RECT 168.860 3.500 174.980 4.300 ;
        RECT 176.140 3.500 182.260 4.300 ;
        RECT 183.420 3.500 189.540 4.300 ;
        RECT 190.700 3.500 196.820 4.300 ;
        RECT 197.980 3.500 204.100 4.300 ;
        RECT 205.260 3.500 211.380 4.300 ;
        RECT 212.540 3.500 218.660 4.300 ;
        RECT 219.820 3.500 225.940 4.300 ;
        RECT 227.100 3.500 233.220 4.300 ;
        RECT 234.380 3.500 240.500 4.300 ;
        RECT 241.660 3.500 247.780 4.300 ;
        RECT 248.940 3.500 255.060 4.300 ;
        RECT 256.220 3.500 262.340 4.300 ;
        RECT 263.500 3.500 269.620 4.300 ;
        RECT 270.780 3.500 276.900 4.300 ;
        RECT 278.060 3.500 284.180 4.300 ;
        RECT 285.340 3.500 291.460 4.300 ;
        RECT 292.620 3.500 298.740 4.300 ;
        RECT 299.900 3.500 306.020 4.300 ;
        RECT 307.180 3.500 313.300 4.300 ;
        RECT 314.460 3.500 320.580 4.300 ;
        RECT 321.740 3.500 327.860 4.300 ;
        RECT 329.020 3.500 335.140 4.300 ;
        RECT 336.300 3.500 342.420 4.300 ;
        RECT 343.580 3.500 349.700 4.300 ;
        RECT 350.860 3.500 356.980 4.300 ;
        RECT 358.140 3.500 364.260 4.300 ;
        RECT 365.420 3.500 371.540 4.300 ;
        RECT 372.700 3.500 378.820 4.300 ;
        RECT 379.980 3.500 386.100 4.300 ;
        RECT 387.260 3.500 393.380 4.300 ;
        RECT 394.540 3.500 400.660 4.300 ;
        RECT 401.820 3.500 407.940 4.300 ;
        RECT 409.100 3.500 415.220 4.300 ;
        RECT 416.380 3.500 422.500 4.300 ;
        RECT 423.660 3.500 429.780 4.300 ;
        RECT 430.940 3.500 437.060 4.300 ;
        RECT 438.220 3.500 444.340 4.300 ;
        RECT 445.500 3.500 451.620 4.300 ;
        RECT 452.780 3.500 458.900 4.300 ;
        RECT 460.060 3.500 466.180 4.300 ;
        RECT 467.340 3.500 473.460 4.300 ;
        RECT 474.620 3.500 480.740 4.300 ;
        RECT 481.900 3.500 488.020 4.300 ;
        RECT 489.180 3.500 495.300 4.300 ;
        RECT 496.460 3.500 502.580 4.300 ;
        RECT 503.740 3.500 509.860 4.300 ;
        RECT 511.020 3.500 517.140 4.300 ;
        RECT 518.300 3.500 524.420 4.300 ;
        RECT 525.580 3.500 531.700 4.300 ;
        RECT 532.860 3.500 538.980 4.300 ;
        RECT 540.140 3.500 546.260 4.300 ;
        RECT 547.420 3.500 553.540 4.300 ;
        RECT 554.700 3.500 560.820 4.300 ;
        RECT 561.980 3.500 568.100 4.300 ;
        RECT 569.260 3.500 575.380 4.300 ;
        RECT 576.540 3.500 582.660 4.300 ;
        RECT 583.820 3.500 589.940 4.300 ;
        RECT 591.100 3.500 597.220 4.300 ;
        RECT 598.380 3.500 604.500 4.300 ;
        RECT 605.660 3.500 611.780 4.300 ;
        RECT 612.940 3.500 619.060 4.300 ;
        RECT 620.220 3.500 626.340 4.300 ;
        RECT 627.500 3.500 633.620 4.300 ;
        RECT 634.780 3.500 640.900 4.300 ;
        RECT 642.060 3.500 648.180 4.300 ;
        RECT 649.340 3.500 655.460 4.300 ;
        RECT 656.620 3.500 662.740 4.300 ;
        RECT 663.900 3.500 670.020 4.300 ;
        RECT 671.180 3.500 677.300 4.300 ;
        RECT 678.460 3.500 684.580 4.300 ;
        RECT 685.740 3.500 691.860 4.300 ;
        RECT 693.020 3.500 699.140 4.300 ;
        RECT 700.300 3.500 706.420 4.300 ;
        RECT 707.580 3.500 713.700 4.300 ;
        RECT 714.860 3.500 720.980 4.300 ;
        RECT 722.140 3.500 728.260 4.300 ;
        RECT 729.420 3.500 735.540 4.300 ;
        RECT 736.700 3.500 742.820 4.300 ;
        RECT 743.980 3.500 750.100 4.300 ;
        RECT 751.260 3.500 757.380 4.300 ;
        RECT 758.540 3.500 764.660 4.300 ;
        RECT 765.820 3.500 771.940 4.300 ;
        RECT 773.100 3.500 779.220 4.300 ;
        RECT 780.380 3.500 786.500 4.300 ;
        RECT 787.660 3.500 793.780 4.300 ;
        RECT 794.940 3.500 801.060 4.300 ;
        RECT 802.220 3.500 808.340 4.300 ;
        RECT 809.500 3.500 815.620 4.300 ;
        RECT 816.780 3.500 822.900 4.300 ;
        RECT 824.060 3.500 830.180 4.300 ;
        RECT 831.340 3.500 837.460 4.300 ;
        RECT 838.620 3.500 844.740 4.300 ;
        RECT 845.900 3.500 852.020 4.300 ;
        RECT 853.180 3.500 859.300 4.300 ;
        RECT 860.460 3.500 866.580 4.300 ;
        RECT 867.740 3.500 873.860 4.300 ;
        RECT 875.020 3.500 881.140 4.300 ;
        RECT 882.300 3.500 888.420 4.300 ;
        RECT 889.580 3.500 895.700 4.300 ;
        RECT 896.860 3.500 902.980 4.300 ;
        RECT 904.140 3.500 910.260 4.300 ;
        RECT 911.420 3.500 917.540 4.300 ;
        RECT 918.700 3.500 924.820 4.300 ;
        RECT 925.980 3.500 932.100 4.300 ;
        RECT 933.260 3.500 939.380 4.300 ;
        RECT 940.540 3.500 946.660 4.300 ;
        RECT 947.820 3.500 953.940 4.300 ;
        RECT 955.100 3.500 961.220 4.300 ;
        RECT 962.380 3.500 968.500 4.300 ;
        RECT 969.660 3.500 975.780 4.300 ;
        RECT 976.940 3.500 983.060 4.300 ;
        RECT 984.220 3.500 990.340 4.300 ;
        RECT 991.500 3.500 991.620 4.300 ;
      LAYER Metal3 ;
        RECT 10.730 14.700 991.670 999.460 ;
      LAYER Metal4 ;
        RECT 515.900 984.520 784.420 998.950 ;
        RECT 515.900 22.490 559.540 984.520 ;
        RECT 561.740 22.490 636.340 984.520 ;
        RECT 638.540 22.490 713.140 984.520 ;
        RECT 715.340 22.490 784.420 984.520 ;
  END
END io_interface
END LIBRARY

