// This is the unpowered netlist.
module io_interface (clk,
    dataw_en,
    hlt,
    instrw_en,
    reset,
    start,
    uP_dataw_en,
    wb_clk_i,
    wb_rst_i,
    data_mem_addr,
    data_read_data,
    data_write_data,
    instr,
    instr_mem_addr,
    instr_write_data,
    io_in,
    io_oeb,
    io_out,
    irq,
    la_data_in,
    la_data_out,
    la_oenb,
    uP_data_mem_addr,
    uP_instr,
    uP_instr_mem_addr,
    uP_write_data);
 output clk;
 output dataw_en;
 input hlt;
 output instrw_en;
 output reset;
 output start;
 input uP_dataw_en;
 input wb_clk_i;
 input wb_rst_i;
 output [7:0] data_mem_addr;
 input [15:0] data_read_data;
 output [15:0] data_write_data;
 input [15:0] instr;
 output [12:0] instr_mem_addr;
 output [15:0] instr_write_data;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [2:0] irq;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 input [7:0] uP_data_mem_addr;
 output [15:0] uP_instr;
 input [12:0] uP_instr_mem_addr;
 input [15:0] uP_write_data;

 wire \Data_out0[0].i2 ;
 wire \Data_out0[0].i3 ;
 wire \Data_out0[10].i3 ;
 wire \Data_out0[11].i3 ;
 wire \Data_out0[12].i3 ;
 wire \Data_out0[1].i2 ;
 wire \Data_out0[1].i3 ;
 wire \Data_out0[2].i2 ;
 wire \Data_out0[2].i3 ;
 wire \Data_out0[3].i2 ;
 wire \Data_out0[3].i3 ;
 wire \Data_out0[4].i2 ;
 wire \Data_out0[4].i3 ;
 wire \Data_out0[5].i2 ;
 wire \Data_out0[5].i3 ;
 wire \Data_out0[6].i2 ;
 wire \Data_out0[6].i3 ;
 wire \Data_out0[7].i2 ;
 wire \Data_out0[7].i3 ;
 wire \Data_out0[8].i3 ;
 wire \Data_out0[9].i3 ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire net356;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net357;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net358;
 wire net313;
 wire net314;
 wire net372;
 wire net373;
 wire net374;
 wire net315;
 wire net375;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net316;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net317;
 wire net318;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;

 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _249_ (.I0(_032_),
    .I1(net55),
    .S(_027_),
    .Z(_108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _250_ (.I(_108_),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _251_ (.I0(_052_),
    .I1(net56),
    .S(_027_),
    .Z(_109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _252_ (.I(_109_),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _253_ (.I0(_058_),
    .I1(net57),
    .S(_027_),
    .Z(_110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _254_ (.I(_110_),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _255_ (.I(_026_),
    .Z(_111_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _256_ (.I0(\Data_out0[3].i2 ),
    .I1(net58),
    .S(_111_),
    .Z(_112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _257_ (.I(_112_),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _258_ (.I0(_068_),
    .I1(net59),
    .S(_111_),
    .Z(_113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _259_ (.I(_113_),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _260_ (.I0(\Data_out0[5].i2 ),
    .I1(net60),
    .S(_111_),
    .Z(_114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _261_ (.I(_114_),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _262_ (.I0(\Data_out0[6].i2 ),
    .I1(net61),
    .S(_111_),
    .Z(_115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _263_ (.I(_115_),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _264_ (.I(_025_),
    .Z(_116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _265_ (.I(_116_),
    .Z(_117_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _266_ (.I0(\Data_out0[7].i2 ),
    .I1(net62),
    .S(_117_),
    .Z(_118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _267_ (.I(_118_),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _268_ (.I0(_044_),
    .I1(net64),
    .S(_117_),
    .Z(_119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _269_ (.I(_119_),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _270_ (.I0(_049_),
    .I1(net68),
    .S(_117_),
    .Z(_120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _271_ (.I(_120_),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _272_ (.I(_025_),
    .Z(_121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _273_ (.I(_121_),
    .Z(_122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _274_ (.I(\Data_out0[2].i3 ),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _275_ (.I(_025_),
    .Z(_124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _276_ (.I(_124_),
    .Z(_125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _277_ (.A1(_125_),
    .A2(net69),
    .ZN(_126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _278_ (.A1(_122_),
    .A2(_123_),
    .B(_126_),
    .ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _279_ (.I0(\Data_out0[3].i3 ),
    .I1(net70),
    .S(_117_),
    .Z(_127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _280_ (.I(_127_),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _281_ (.I(_116_),
    .Z(_128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _282_ (.I0(_069_),
    .I1(net71),
    .S(_128_),
    .Z(_129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _283_ (.I(_129_),
    .Z(net128));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _284_ (.I0(\Data_out0[5].i3 ),
    .I1(net72),
    .S(_128_),
    .Z(_130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _285_ (.I(_130_),
    .Z(net129));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _286_ (.I0(_077_),
    .I1(net73),
    .S(_128_),
    .Z(_131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _287_ (.I(_131_),
    .Z(net130));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _288_ (.I0(\Data_out0[7].i3 ),
    .I1(net74),
    .S(_128_),
    .Z(_132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _289_ (.I(_132_),
    .Z(net131));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _290_ (.I(_116_),
    .Z(_133_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _291_ (.I0(_085_),
    .I1(net75),
    .S(_133_),
    .Z(_134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _292_ (.I(_134_),
    .Z(net132));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _293_ (.I0(\Data_out0[9].i3 ),
    .I1(net76),
    .S(_133_),
    .Z(_135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _294_ (.I(_135_),
    .Z(net133));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _295_ (.I0(_093_),
    .I1(net65),
    .S(_133_),
    .Z(_136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _296_ (.I(_136_),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _297_ (.I0(\Data_out0[11].i3 ),
    .I1(net66),
    .S(_133_),
    .Z(_137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _298_ (.I(_137_),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _299_ (.I(_116_),
    .Z(_138_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _300_ (.I0(\Data_out0[12].i3 ),
    .I1(net67),
    .S(_138_),
    .Z(_139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _301_ (.I(_139_),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _302_ (.I(_026_),
    .Z(_140_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _303_ (.A1(_140_),
    .A2(net18),
    .Z(_141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _304_ (.I(_141_),
    .Z(net196));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _305_ (.A1(_140_),
    .A2(net25),
    .Z(_142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _306_ (.I(_142_),
    .Z(net197));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _307_ (.A1(_023_),
    .A2(net26),
    .Z(_143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _308_ (.I(_143_),
    .Z(net198));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _309_ (.A1(_140_),
    .A2(net27),
    .Z(_144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _310_ (.I(_144_),
    .Z(net199));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _311_ (.I(_121_),
    .Z(_145_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _312_ (.A1(_145_),
    .A2(net28),
    .Z(_146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _313_ (.I(_146_),
    .Z(net200));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _314_ (.A1(_145_),
    .A2(net29),
    .Z(_147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _315_ (.I(_147_),
    .Z(net201));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _316_ (.A1(_145_),
    .A2(net30),
    .Z(_148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _317_ (.I(_148_),
    .Z(net202));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _318_ (.A1(_145_),
    .A2(net31),
    .Z(_149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _319_ (.I(_149_),
    .Z(net203));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _320_ (.I(_026_),
    .Z(_150_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _321_ (.A1(_150_),
    .A2(net32),
    .Z(_151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _322_ (.I(_151_),
    .Z(net204));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _323_ (.A1(_150_),
    .A2(net33),
    .Z(_152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _324_ (.I(_152_),
    .Z(net205));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _325_ (.A1(_150_),
    .A2(net19),
    .Z(_153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _326_ (.I(_153_),
    .Z(net206));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _327_ (.A1(_150_),
    .A2(net20),
    .Z(_154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _328_ (.I(_154_),
    .Z(net207));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _329_ (.A1(_125_),
    .A2(net21),
    .Z(_155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _330_ (.I(_155_),
    .Z(net208));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _331_ (.A1(_023_),
    .A2(net22),
    .Z(_156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _332_ (.I(_156_),
    .Z(net209));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _333_ (.A1(_125_),
    .A2(net23),
    .Z(_157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _334_ (.I(_157_),
    .Z(net210));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _335_ (.A1(_125_),
    .A2(net24),
    .Z(_158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _336_ (.I(_158_),
    .Z(net211));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _337_ (.I(net63),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _338_ (.A1(_021_),
    .A2(_034_),
    .A3(_024_),
    .B1(_159_),
    .B2(_023_),
    .ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _339_ (.I(_124_),
    .Z(_160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _340_ (.A1(_160_),
    .A2(net77),
    .ZN(_161_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _341_ (.A1(_122_),
    .A2(_029_),
    .B(_161_),
    .ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _342_ (.A1(_160_),
    .A2(net84),
    .ZN(_162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _343_ (.A1(_122_),
    .A2(_048_),
    .B(_162_),
    .ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _344_ (.A1(_160_),
    .A2(net85),
    .ZN(_163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _345_ (.A1(_122_),
    .A2(_055_),
    .B(_163_),
    .ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _346_ (.I(_121_),
    .Z(_164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _347_ (.A1(_160_),
    .A2(net86),
    .ZN(_165_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _348_ (.A1(_164_),
    .A2(_061_),
    .B(_165_),
    .ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _349_ (.I(_124_),
    .Z(_166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _350_ (.A1(_166_),
    .A2(net87),
    .ZN(_167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _351_ (.A1(_164_),
    .A2(_065_),
    .B(_167_),
    .ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _352_ (.A1(_166_),
    .A2(net88),
    .ZN(_168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _353_ (.A1(_164_),
    .A2(_071_),
    .B(_168_),
    .ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _354_ (.A1(_166_),
    .A2(net89),
    .ZN(_169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _355_ (.A1(_164_),
    .A2(_076_),
    .B(_169_),
    .ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _356_ (.A1(_166_),
    .A2(net90),
    .ZN(_170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _357_ (.A1(_140_),
    .A2(_080_),
    .B(_170_),
    .ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _358_ (.I0(net53),
    .I1(net91),
    .S(_138_),
    .Z(_171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _359_ (.I(_171_),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _360_ (.I0(net54),
    .I1(net92),
    .S(_138_),
    .Z(_172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _361_ (.I(_172_),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _362_ (.I0(net35),
    .I1(net78),
    .S(_138_),
    .Z(_173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _363_ (.I(_173_),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _364_ (.I(_124_),
    .Z(_174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _365_ (.I0(net36),
    .I1(net79),
    .S(_174_),
    .Z(_175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _366_ (.I(_175_),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _367_ (.I0(net37),
    .I1(net80),
    .S(_174_),
    .Z(_176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _368_ (.I(_176_),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _369_ (.I0(net38),
    .I1(net81),
    .S(_174_),
    .Z(_177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _370_ (.I(_177_),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _371_ (.I0(net39),
    .I1(net82),
    .S(_174_),
    .Z(_178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _372_ (.I(_178_),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _373_ (.I0(net40),
    .I1(net83),
    .S(_121_),
    .Z(_179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _374_ (.I(_179_),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _375_ (.A1(_033_),
    .A2(_034_),
    .A3(_024_),
    .ZN(_180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _376_ (.I(_180_),
    .Z(_181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _377_ (.I(_180_),
    .Z(_182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _378_ (.A1(net34),
    .A2(_182_),
    .ZN(_183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _379_ (.A1(_032_),
    .A2(_181_),
    .B(_183_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _380_ (.A1(\Data_out0[0].i2 ),
    .A2(\Data_out0[1].i2 ),
    .ZN(_184_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _381_ (.A1(_032_),
    .A2(_052_),
    .Z(_185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _382_ (.I(_180_),
    .Z(_186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _383_ (.A1(_184_),
    .A2(_185_),
    .B(_186_),
    .ZN(_187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _384_ (.A1(_048_),
    .A2(_181_),
    .B(_187_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _385_ (.I(_180_),
    .Z(_188_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _386_ (.A1(_058_),
    .A2(_184_),
    .Z(_189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _387_ (.A1(net42),
    .A2(_182_),
    .ZN(_190_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _388_ (.A1(_188_),
    .A2(_189_),
    .B(_190_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _389_ (.A1(\Data_out0[0].i2 ),
    .A2(_052_),
    .A3(_058_),
    .ZN(_191_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _390_ (.A1(\Data_out0[3].i2 ),
    .A2(_191_),
    .Z(_192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _391_ (.A1(net48),
    .A2(_182_),
    .ZN(_193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _392_ (.A1(_188_),
    .A2(_192_),
    .B(_193_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _393_ (.A1(\Data_out0[0].i2 ),
    .A2(\Data_out0[1].i2 ),
    .A3(\Data_out0[2].i2 ),
    .A4(\Data_out0[3].i2 ),
    .Z(_194_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _394_ (.A1(_068_),
    .A2(_194_),
    .Z(_195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _395_ (.A1(_186_),
    .A2(_195_),
    .ZN(_196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _396_ (.A1(_065_),
    .A2(_181_),
    .B(_196_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _397_ (.A1(_068_),
    .A2(_194_),
    .B(\Data_out0[5].i2 ),
    .ZN(_197_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _398_ (.A1(\Data_out0[4].i2 ),
    .A2(\Data_out0[5].i2 ),
    .A3(_194_),
    .Z(_198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _399_ (.A1(net50),
    .A2(_186_),
    .ZN(_199_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _400_ (.A1(_188_),
    .A2(_197_),
    .A3(_198_),
    .B(_199_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _401_ (.A1(\Data_out0[6].i2 ),
    .A2(_198_),
    .Z(_200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _402_ (.A1(\Data_out0[6].i2 ),
    .A2(_198_),
    .ZN(_201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _403_ (.A1(_200_),
    .A2(_201_),
    .B(_186_),
    .ZN(_202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _404_ (.A1(_076_),
    .A2(_181_),
    .B(_202_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _405_ (.A1(\Data_out0[7].i2 ),
    .A2(_201_),
    .Z(_203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _406_ (.A1(net52),
    .A2(_182_),
    .ZN(_204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _407_ (.A1(_188_),
    .A2(_203_),
    .B(_204_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _408_ (.A1(_033_),
    .A2(_022_),
    .A3(_024_),
    .ZN(_205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _409_ (.I(_205_),
    .Z(_206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _410_ (.I(_206_),
    .Z(_207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _411_ (.I(_205_),
    .Z(_208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _412_ (.A1(net34),
    .A2(_208_),
    .ZN(_209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _413_ (.A1(_044_),
    .A2(_207_),
    .B(_209_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _414_ (.I(_206_),
    .Z(_210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _415_ (.A1(\Data_out0[0].i3 ),
    .A2(_049_),
    .ZN(_211_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _416_ (.A1(_044_),
    .A2(_049_),
    .Z(_212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _417_ (.I(_205_),
    .Z(_213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _418_ (.A1(_211_),
    .A2(_212_),
    .B(_213_),
    .ZN(_214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _419_ (.A1(_048_),
    .A2(_210_),
    .B(_214_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _420_ (.A1(\Data_out0[0].i3 ),
    .A2(\Data_out0[1].i3 ),
    .A3(\Data_out0[2].i3 ),
    .ZN(_215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _421_ (.A1(_123_),
    .A2(_211_),
    .ZN(_216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _422_ (.A1(_215_),
    .A2(_216_),
    .B(_206_),
    .ZN(_217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _423_ (.A1(_055_),
    .A2(_210_),
    .B(_217_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _424_ (.A1(\Data_out0[3].i3 ),
    .A2(_215_),
    .Z(_218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _425_ (.A1(net48),
    .A2(_208_),
    .ZN(_219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _426_ (.A1(_207_),
    .A2(_218_),
    .B(_219_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _427_ (.A1(\Data_out0[0].i3 ),
    .A2(\Data_out0[1].i3 ),
    .A3(\Data_out0[2].i3 ),
    .A4(\Data_out0[3].i3 ),
    .Z(_220_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _428_ (.A1(_069_),
    .A2(_220_),
    .Z(_221_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _429_ (.A1(_213_),
    .A2(_221_),
    .ZN(_222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _430_ (.A1(_065_),
    .A2(_210_),
    .B(_222_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _431_ (.I(_206_),
    .Z(_223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _432_ (.A1(_069_),
    .A2(_220_),
    .B(\Data_out0[5].i3 ),
    .ZN(_224_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _433_ (.A1(\Data_out0[4].i3 ),
    .A2(\Data_out0[5].i3 ),
    .Z(_225_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _434_ (.A1(_220_),
    .A2(_225_),
    .Z(_226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _435_ (.I(_205_),
    .Z(_227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _436_ (.A1(net50),
    .A2(_227_),
    .ZN(_228_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _437_ (.A1(_223_),
    .A2(_224_),
    .A3(_226_),
    .B(_228_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _438_ (.A1(_077_),
    .A2(_226_),
    .Z(_229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _439_ (.A1(_213_),
    .A2(_229_),
    .ZN(_230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _440_ (.A1(_076_),
    .A2(_210_),
    .B(_230_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _441_ (.A1(_077_),
    .A2(_226_),
    .B(\Data_out0[7].i3 ),
    .ZN(_231_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _442_ (.A1(\Data_out0[6].i3 ),
    .A2(\Data_out0[7].i3 ),
    .A3(_220_),
    .A4(_225_),
    .Z(_232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _443_ (.I(_232_),
    .Z(_233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _444_ (.A1(net52),
    .A2(_227_),
    .ZN(_234_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _445_ (.A1(_223_),
    .A2(_231_),
    .A3(_233_),
    .B(_234_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _446_ (.A1(_085_),
    .A2(_233_),
    .Z(_235_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _447_ (.I0(_235_),
    .I1(net53),
    .S(_213_),
    .Z(_236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _448_ (.I(_236_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _449_ (.A1(_085_),
    .A2(_233_),
    .B(\Data_out0[9].i3 ),
    .ZN(_237_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _450_ (.A1(\Data_out0[8].i3 ),
    .A2(\Data_out0[9].i3 ),
    .Z(_238_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _451_ (.A1(_232_),
    .A2(_238_),
    .Z(_239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _452_ (.A1(net54),
    .A2(_227_),
    .ZN(_240_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _453_ (.A1(_223_),
    .A2(_237_),
    .A3(_239_),
    .B(_240_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _454_ (.A1(_093_),
    .A2(_239_),
    .ZN(_241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _455_ (.A1(net35),
    .A2(_208_),
    .ZN(_242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _456_ (.A1(_207_),
    .A2(_241_),
    .B(_242_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _457_ (.A1(_093_),
    .A2(_233_),
    .A3(_238_),
    .ZN(_243_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _458_ (.A1(\Data_out0[11].i3 ),
    .A2(_243_),
    .Z(_244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _459_ (.A1(net36),
    .A2(_208_),
    .ZN(_245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _460_ (.A1(_207_),
    .A2(_244_),
    .B(_245_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _461_ (.A1(\Data_out0[10].i3 ),
    .A2(\Data_out0[11].i3 ),
    .A3(_232_),
    .A4(_238_),
    .ZN(_246_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _462_ (.A1(\Data_out0[12].i3 ),
    .A2(_246_),
    .Z(_247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _463_ (.A1(net37),
    .A2(_227_),
    .ZN(_248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _464_ (.A1(_223_),
    .A2(_247_),
    .B(_248_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _465_ (.I(net45),
    .Z(_021_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _466_ (.I(net44),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _467_ (.I(net46),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _468_ (.A1(_023_),
    .A2(net43),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _469_ (.A1(_021_),
    .A2(_022_),
    .A3(_024_),
    .ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _470_ (.I(net46),
    .Z(_025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _471_ (.I(_025_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _472_ (.I(_026_),
    .Z(_027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _473_ (.I0(net47),
    .I1(net93),
    .S(_027_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _474_ (.I(_028_),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _475_ (.I(net34),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _476_ (.I(net43),
    .Z(_030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _477_ (.I(_030_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _478_ (.I(\Data_out0[0].i2 ),
    .Z(_032_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _479_ (.I(net45),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _480_ (.I(net44),
    .Z(_034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _481_ (.A1(_033_),
    .A2(_034_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _482_ (.I(_035_),
    .Z(_036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _483_ (.I(net43),
    .Z(_037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _484_ (.I(_037_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _485_ (.A1(_032_),
    .A2(_036_),
    .B(_038_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _486_ (.A1(_021_),
    .A2(_022_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _487_ (.I(_040_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _488_ (.A1(_033_),
    .A2(_022_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _489_ (.I(_042_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _490_ (.I(\Data_out0[0].i3 ),
    .Z(_044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _491_ (.A1(_021_),
    .A2(_034_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _492_ (.I(_045_),
    .Z(_046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _493_ (.A1(net18),
    .A2(_041_),
    .B1(_043_),
    .B2(_044_),
    .C1(_046_),
    .C2(net1),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _494_ (.A1(_029_),
    .A2(_031_),
    .B1(_039_),
    .B2(_047_),
    .ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _495_ (.I(net41),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _496_ (.I(\Data_out0[1].i3 ),
    .Z(_049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _497_ (.A1(_049_),
    .A2(_043_),
    .B(_038_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _498_ (.I(_035_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _499_ (.I(\Data_out0[1].i2 ),
    .Z(_052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _500_ (.I(_045_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _501_ (.A1(net25),
    .A2(_041_),
    .B1(_051_),
    .B2(_052_),
    .C1(_053_),
    .C2(net8),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _502_ (.A1(_031_),
    .A2(_048_),
    .B1(_050_),
    .B2(_054_),
    .ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _503_ (.I(net42),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _504_ (.I(_040_),
    .Z(_056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _505_ (.A1(net26),
    .A2(_056_),
    .B(_038_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _506_ (.I(\Data_out0[2].i2 ),
    .Z(_058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _507_ (.I(_042_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _508_ (.A1(_058_),
    .A2(_036_),
    .B1(_059_),
    .B2(\Data_out0[2].i3 ),
    .C1(_053_),
    .C2(net9),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _509_ (.A1(_031_),
    .A2(_055_),
    .B1(_057_),
    .B2(_060_),
    .ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _510_ (.I(net48),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _511_ (.A1(\Data_out0[3].i3 ),
    .A2(_043_),
    .B(_038_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _512_ (.A1(net27),
    .A2(_041_),
    .B1(_051_),
    .B2(\Data_out0[3].i2 ),
    .C1(_053_),
    .C2(net10),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _513_ (.A1(_031_),
    .A2(_061_),
    .B1(_062_),
    .B2(_063_),
    .ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _514_ (.I(_030_),
    .Z(_064_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _515_ (.I(net49),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _516_ (.I(_037_),
    .Z(_066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _517_ (.A1(net28),
    .A2(_056_),
    .B(_066_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _518_ (.I(\Data_out0[4].i2 ),
    .Z(_068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _519_ (.I(\Data_out0[4].i3 ),
    .Z(_069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _520_ (.A1(_068_),
    .A2(_051_),
    .B1(_059_),
    .B2(_069_),
    .C1(_053_),
    .C2(net11),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _521_ (.A1(_064_),
    .A2(_065_),
    .B1(_067_),
    .B2(_070_),
    .ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _522_ (.I(net50),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _523_ (.A1(\Data_out0[5].i2 ),
    .A2(_036_),
    .B(_066_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _524_ (.I(_040_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _525_ (.I(_045_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _526_ (.A1(net29),
    .A2(_073_),
    .B1(_059_),
    .B2(\Data_out0[5].i3 ),
    .C1(_074_),
    .C2(net12),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _527_ (.A1(_064_),
    .A2(_071_),
    .B1(_072_),
    .B2(_075_),
    .ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _528_ (.I(net51),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _529_ (.I(\Data_out0[6].i3 ),
    .Z(_077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _530_ (.A1(_077_),
    .A2(_043_),
    .B(_066_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _531_ (.A1(net30),
    .A2(_073_),
    .B1(_051_),
    .B2(\Data_out0[6].i2 ),
    .C1(_074_),
    .C2(net13),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _532_ (.A1(_064_),
    .A2(_076_),
    .B1(_078_),
    .B2(_079_),
    .ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _533_ (.I(net52),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _534_ (.A1(\Data_out0[7].i2 ),
    .A2(_036_),
    .B(_066_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _535_ (.A1(net31),
    .A2(_073_),
    .B1(_059_),
    .B2(\Data_out0[7].i3 ),
    .C1(_074_),
    .C2(net14),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _536_ (.A1(_064_),
    .A2(_080_),
    .B1(_081_),
    .B2(_082_),
    .ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _537_ (.I(_030_),
    .Z(_083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _538_ (.I(_042_),
    .Z(_084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _539_ (.I(\Data_out0[8].i3 ),
    .Z(_085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _540_ (.A1(net32),
    .A2(_073_),
    .B1(_084_),
    .B2(_085_),
    .C1(_074_),
    .C2(net15),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _541_ (.I(_037_),
    .Z(_087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _542_ (.A1(_087_),
    .A2(net53),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _543_ (.A1(_083_),
    .A2(_086_),
    .B(_088_),
    .ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _544_ (.I(_040_),
    .Z(_089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _545_ (.I(_045_),
    .Z(_090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _546_ (.A1(net33),
    .A2(_089_),
    .B1(_084_),
    .B2(\Data_out0[9].i3 ),
    .C1(_090_),
    .C2(net16),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _547_ (.A1(_087_),
    .A2(net54),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _548_ (.A1(_083_),
    .A2(_091_),
    .B(_092_),
    .ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _549_ (.I(\Data_out0[10].i3 ),
    .Z(_093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _550_ (.A1(net19),
    .A2(_089_),
    .B1(_084_),
    .B2(_093_),
    .C1(_090_),
    .C2(net2),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _551_ (.A1(_087_),
    .A2(net35),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _552_ (.A1(_083_),
    .A2(_094_),
    .B(_095_),
    .ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _553_ (.A1(net20),
    .A2(_089_),
    .B1(_084_),
    .B2(\Data_out0[11].i3 ),
    .C1(_090_),
    .C2(net3),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _554_ (.A1(_087_),
    .A2(net36),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _555_ (.A1(_083_),
    .A2(_096_),
    .B(_097_),
    .ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _556_ (.I(_030_),
    .Z(_098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _557_ (.A1(net21),
    .A2(_089_),
    .B1(_042_),
    .B2(\Data_out0[12].i3 ),
    .C1(_090_),
    .C2(net4),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _558_ (.I(_037_),
    .Z(_100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _559_ (.A1(_100_),
    .A2(net37),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _560_ (.A1(_098_),
    .A2(_099_),
    .B(_101_),
    .ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _561_ (.A1(net22),
    .A2(_056_),
    .B1(_046_),
    .B2(net5),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _562_ (.A1(_100_),
    .A2(net38),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _563_ (.A1(_098_),
    .A2(_102_),
    .B(_103_),
    .ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _564_ (.A1(net23),
    .A2(_056_),
    .B1(_046_),
    .B2(net6),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _565_ (.A1(_100_),
    .A2(net39),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _566_ (.A1(_098_),
    .A2(_104_),
    .B(_105_),
    .ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _567_ (.A1(net24),
    .A2(_041_),
    .B1(_046_),
    .B2(net7),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _568_ (.A1(_100_),
    .A2(net40),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _569_ (.A1(_098_),
    .A2(_106_),
    .B(_107_),
    .ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _570_ (.D(_000_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[0].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _571_ (.D(_001_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[1].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _572_ (.D(_002_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[2].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _573_ (.D(_003_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[3].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _574_ (.D(_004_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[4].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _575_ (.D(_005_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[5].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _576_ (.D(_006_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[6].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _577_ (.D(_007_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[7].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _578_ (.D(_008_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[0].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _579_ (.D(_012_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[1].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _580_ (.D(_013_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[2].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _581_ (.D(_014_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[3].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _582_ (.D(_015_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[4].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _583_ (.D(_016_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[5].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _584_ (.D(_017_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[6].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _585_ (.D(_018_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[7].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _586_ (.D(_019_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[8].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _587_ (.D(_020_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[9].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _588_ (.D(_009_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[10].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _589_ (.D(_010_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[11].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _590_ (.D(_011_),
    .RN(net94),
    .CLK(net95),
    .Q(\Data_out0[12].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_356 (.Z(net356));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_357 (.Z(net357));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_358 (.Z(net358));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_359 (.Z(net359));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_360 (.Z(net360));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_361 (.Z(net361));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_362 (.Z(net362));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_363 (.Z(net363));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_364 (.Z(net364));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_365 (.Z(net365));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_366 (.Z(net366));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_367 (.Z(net367));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_368 (.Z(net368));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_369 (.Z(net369));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_370 (.Z(net370));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_371 (.Z(net371));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_372 (.Z(net372));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_373 (.Z(net373));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_374 (.Z(net374));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_375 (.Z(net375));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__553__B2 (.I(\Data_out0[11].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_299 (.ZN(net299));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_300 (.ZN(net300));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_301 (.ZN(net301));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_302 (.ZN(net302));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_303 (.ZN(net303));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_304 (.ZN(net304));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_305 (.ZN(net305));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_306 (.ZN(net306));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_307 (.ZN(net307));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_308 (.ZN(net308));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_309 (.ZN(net309));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_310 (.ZN(net310));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_311 (.ZN(net311));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_312 (.ZN(net312));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_313 (.ZN(net313));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_314 (.ZN(net314));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_315 (.ZN(net315));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_316 (.ZN(net316));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_317 (.ZN(net317));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_318 (.ZN(net318));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_319 (.ZN(net319));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_320 (.ZN(net320));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_321 (.ZN(net321));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_322 (.ZN(net322));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_323 (.ZN(net323));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_324 (.ZN(net324));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_325 (.ZN(net325));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_326 (.ZN(net326));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_327 (.ZN(net327));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_328 (.ZN(net328));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_329 (.ZN(net329));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_330 (.ZN(net330));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_331 (.ZN(net331));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_332 (.ZN(net332));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_333 (.ZN(net333));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_334 (.ZN(net334));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_335 (.ZN(net335));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_336 (.ZN(net336));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_337 (.ZN(net337));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_338 (.ZN(net338));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_339 (.ZN(net339));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_340 (.ZN(net340));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_341 (.ZN(net341));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_342 (.ZN(net342));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_343 (.ZN(net343));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_344 (.ZN(net344));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_345 (.ZN(net345));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_346 (.ZN(net346));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_347 (.ZN(net347));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_348 (.ZN(net348));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_349 (.ZN(net349));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_350 (.ZN(net350));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_351 (.ZN(net351));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_352 (.ZN(net352));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_353 (.ZN(net353));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_354 (.ZN(net354));
 gf180mcu_fd_sc_mcu7t5v0__tieh io_interface_355 (.Z(net355));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _669_ (.I(net34),
    .Z(net134));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _670_ (.I(net41),
    .Z(net141));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _671_ (.I(net42),
    .Z(net142));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _672_ (.I(net48),
    .Z(net143));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _673_ (.I(net49),
    .Z(net144));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _674_ (.I(net50),
    .Z(net145));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _675_ (.I(net51),
    .Z(net146));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _676_ (.I(net52),
    .Z(net147));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _677_ (.I(net53),
    .Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _678_ (.I(net54),
    .Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _679_ (.I(net35),
    .Z(net135));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _680_ (.I(net36),
    .Z(net136));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _681_ (.I(net37),
    .Z(net137));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _682_ (.I(net38),
    .Z(net138));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _683_ (.I(net39),
    .Z(net139));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _684_ (.I(net40),
    .Z(net140));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _685_ (.I(net17),
    .Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _686_ (.I(net121),
    .Z(net212));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _687_ (.I(net125),
    .Z(net213));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _688_ (.I(net126),
    .Z(net214));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _689_ (.I(net127),
    .Z(net215));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _690_ (.I(net128),
    .Z(net216));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _691_ (.I(net129),
    .Z(net217));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _692_ (.I(net130),
    .Z(net218));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _693_ (.I(net131),
    .Z(net219));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _694_ (.I(net132),
    .Z(net220));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _695_ (.I(net133),
    .Z(net221));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _696_ (.I(net122),
    .Z(net222));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _697_ (.I(net123),
    .Z(net223));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _698_ (.I(net124),
    .Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _699_ (.I(net104),
    .Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _700_ (.I(net111),
    .Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _701_ (.I(net112),
    .Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _702_ (.I(net113),
    .Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _703_ (.I(net114),
    .Z(net229));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _704_ (.I(net115),
    .Z(net230));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _705_ (.I(net116),
    .Z(net231));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _706_ (.I(net117),
    .Z(net232));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _707_ (.I(net118),
    .Z(net233));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _708_ (.I(net119),
    .Z(net234));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _709_ (.I(net105),
    .Z(net235));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _710_ (.I(net106),
    .Z(net236));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _711_ (.I(net107),
    .Z(net237));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _712_ (.I(net108),
    .Z(net238));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _713_ (.I(net109),
    .Z(net239));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _714_ (.I(net110),
    .Z(net240));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _715_ (.I(net1),
    .Z(net241));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _716_ (.I(net8),
    .Z(net242));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _717_ (.I(net9),
    .Z(net243));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _718_ (.I(net10),
    .Z(net244));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _719_ (.I(net11),
    .Z(net245));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _720_ (.I(net12),
    .Z(net246));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _721_ (.I(net13),
    .Z(net247));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _722_ (.I(net14),
    .Z(net248));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _723_ (.I(net15),
    .Z(net249));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _724_ (.I(net16),
    .Z(net250));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _725_ (.I(net2),
    .Z(net251));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _726_ (.I(net3),
    .Z(net252));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _727_ (.I(net4),
    .Z(net253));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _728_ (.I(net5),
    .Z(net254));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _729_ (.I(net6),
    .Z(net255));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _730_ (.I(net7),
    .Z(net256));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _731_ (.I(net96),
    .Z(net257));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _732_ (.I(net97),
    .Z(net258));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _733_ (.I(net98),
    .Z(net259));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _734_ (.I(net99),
    .Z(net260));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _735_ (.I(net100),
    .Z(net261));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _736_ (.I(net101),
    .Z(net262));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _737_ (.I(net102),
    .Z(net263));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _738_ (.I(net103),
    .Z(net264));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _739_ (.I(net151),
    .Z(net265));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _740_ (.I(net152),
    .Z(net266));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _741_ (.I(net153),
    .Z(net267));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _742_ (.I(net154),
    .Z(net268));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _743_ (.I(net155),
    .Z(net269));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _744_ (.I(net156),
    .Z(net270));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _745_ (.I(net157),
    .Z(net271));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _746_ (.I(net158),
    .Z(net272));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _747_ (.I(net159),
    .Z(net273));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _748_ (.I(net160),
    .Z(net274));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _749_ (.I(net161),
    .Z(net275));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _750_ (.I(net162),
    .Z(net276));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _751_ (.I(net163),
    .Z(net277));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _752_ (.I(net164),
    .Z(net278));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _753_ (.I(net165),
    .Z(net279));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _754_ (.I(net166),
    .Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _755_ (.I(net43),
    .Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _756_ (.I(net44),
    .Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _757_ (.I(net45),
    .Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _758_ (.I(net34),
    .Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _759_ (.I(net41),
    .Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _760_ (.I(net42),
    .Z(net174));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _761_ (.I(net48),
    .Z(net175));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _762_ (.I(net49),
    .Z(net176));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _763_ (.I(net50),
    .Z(net177));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _764_ (.I(net51),
    .Z(net178));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _765_ (.I(net52),
    .Z(net179));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _766_ (.I(net53),
    .Z(net180));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _767_ (.I(net54),
    .Z(net181));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _768_ (.I(net35),
    .Z(net182));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _769_ (.I(net36),
    .Z(net183));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _770_ (.I(net37),
    .Z(net184));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _771_ (.I(net38),
    .Z(net185));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _772_ (.I(net39),
    .Z(net186));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _773_ (.I(net40),
    .Z(net187));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _774_ (.I(net46),
    .Z(net188));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _775_ (.I(net150),
    .Z(net189));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _776_ (.I(net120),
    .Z(net190));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _777_ (.I(net63),
    .Z(net191));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _778_ (.I(net94),
    .Z(net192));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _779_ (.I(net47),
    .Z(net193));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _780_ (.I(net93),
    .Z(net194));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _781_ (.I(net95),
    .Z(net195));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _782_ (.I(net94),
    .Z(net280));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _783_ (.I(net46),
    .Z(net281));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _784_ (.I(net196),
    .Z(net282));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _785_ (.I(net197),
    .Z(net289));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _786_ (.I(net198),
    .Z(net290));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _787_ (.I(net199),
    .Z(net291));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _788_ (.I(net200),
    .Z(net292));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _789_ (.I(net201),
    .Z(net293));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _790_ (.I(net202),
    .Z(net294));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _791_ (.I(net203),
    .Z(net295));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _792_ (.I(net204),
    .Z(net296));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _793_ (.I(net205),
    .Z(net297));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _794_ (.I(net206),
    .Z(net283));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _795_ (.I(net207),
    .Z(net284));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _796_ (.I(net208),
    .Z(net285));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _797_ (.I(net209),
    .Z(net286));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _798_ (.I(net210),
    .Z(net287));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _799_ (.I(net211),
    .Z(net288));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(data_read_data[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(data_read_data[10]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(data_read_data[11]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(data_read_data[12]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(data_read_data[13]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(data_read_data[14]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(data_read_data[15]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(data_read_data[1]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(data_read_data[2]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(data_read_data[3]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(data_read_data[4]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(data_read_data[5]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(data_read_data[6]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(data_read_data[7]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(data_read_data[8]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(data_read_data[9]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(hlt),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(instr[0]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(instr[10]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(instr[11]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(instr[12]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(instr[13]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(instr[14]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(instr[15]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(instr[1]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(instr[2]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(instr[3]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(instr[4]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(instr[5]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(instr[6]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(instr[7]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(instr[8]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(instr[9]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input34 (.I(io_in[0]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input35 (.I(io_in[10]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input36 (.I(io_in[11]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input37 (.I(io_in[12]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input38 (.I(io_in[13]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input39 (.I(io_in[14]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input40 (.I(io_in[15]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input41 (.I(io_in[1]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input42 (.I(io_in[2]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input43 (.I(io_in[32]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input44 (.I(io_in[33]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input45 (.I(io_in[34]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input46 (.I(io_in[36]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input47 (.I(io_in[37]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input48 (.I(io_in[3]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input49 (.I(io_in[4]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input50 (.I(io_in[5]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input51 (.I(io_in[6]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input52 (.I(io_in[7]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input53 (.I(io_in[8]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input54 (.I(io_in[9]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input55 (.I(uP_data_mem_addr[0]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input56 (.I(uP_data_mem_addr[1]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input57 (.I(uP_data_mem_addr[2]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input58 (.I(uP_data_mem_addr[3]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input59 (.I(uP_data_mem_addr[4]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input60 (.I(uP_data_mem_addr[5]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input61 (.I(uP_data_mem_addr[6]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input62 (.I(uP_data_mem_addr[7]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input63 (.I(uP_dataw_en),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input64 (.I(uP_instr_mem_addr[0]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input65 (.I(uP_instr_mem_addr[10]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input66 (.I(uP_instr_mem_addr[11]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input67 (.I(uP_instr_mem_addr[12]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input68 (.I(uP_instr_mem_addr[1]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input69 (.I(uP_instr_mem_addr[2]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input70 (.I(uP_instr_mem_addr[3]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input71 (.I(uP_instr_mem_addr[4]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input72 (.I(uP_instr_mem_addr[5]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input73 (.I(uP_instr_mem_addr[6]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input74 (.I(uP_instr_mem_addr[7]),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input75 (.I(uP_instr_mem_addr[8]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input76 (.I(uP_instr_mem_addr[9]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input77 (.I(uP_write_data[0]),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input78 (.I(uP_write_data[10]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input79 (.I(uP_write_data[11]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input80 (.I(uP_write_data[12]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input81 (.I(uP_write_data[13]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input82 (.I(uP_write_data[14]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input83 (.I(uP_write_data[15]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input84 (.I(uP_write_data[1]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input85 (.I(uP_write_data[2]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input86 (.I(uP_write_data[3]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input87 (.I(uP_write_data[4]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input88 (.I(uP_write_data[5]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input89 (.I(uP_write_data[6]),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input90 (.I(uP_write_data[7]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input91 (.I(uP_write_data[8]),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input92 (.I(uP_write_data[9]),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input93 (.I(wb_clk_i),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input94 (.I(wb_rst_i),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output95 (.I(net95),
    .Z(clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output96 (.I(net96),
    .Z(data_mem_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output97 (.I(net97),
    .Z(data_mem_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output98 (.I(net98),
    .Z(data_mem_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output99 (.I(net99),
    .Z(data_mem_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output100 (.I(net100),
    .Z(data_mem_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output101 (.I(net101),
    .Z(data_mem_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output102 (.I(net102),
    .Z(data_mem_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output103 (.I(net103),
    .Z(data_mem_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output104 (.I(net104),
    .Z(data_write_data[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output105 (.I(net105),
    .Z(data_write_data[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output106 (.I(net106),
    .Z(data_write_data[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output107 (.I(net107),
    .Z(data_write_data[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output108 (.I(net108),
    .Z(data_write_data[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output109 (.I(net109),
    .Z(data_write_data[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output110 (.I(net110),
    .Z(data_write_data[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output111 (.I(net111),
    .Z(data_write_data[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output112 (.I(net112),
    .Z(data_write_data[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output113 (.I(net113),
    .Z(data_write_data[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output114 (.I(net114),
    .Z(data_write_data[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output115 (.I(net115),
    .Z(data_write_data[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output116 (.I(net116),
    .Z(data_write_data[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output117 (.I(net117),
    .Z(data_write_data[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output118 (.I(net118),
    .Z(data_write_data[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output119 (.I(net119),
    .Z(data_write_data[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output120 (.I(net120),
    .Z(dataw_en));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output121 (.I(net121),
    .Z(instr_mem_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output122 (.I(net122),
    .Z(instr_mem_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output123 (.I(net123),
    .Z(instr_mem_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output124 (.I(net124),
    .Z(instr_mem_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output125 (.I(net125),
    .Z(instr_mem_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output126 (.I(net126),
    .Z(instr_mem_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output127 (.I(net127),
    .Z(instr_mem_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output128 (.I(net128),
    .Z(instr_mem_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output129 (.I(net129),
    .Z(instr_mem_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output130 (.I(net130),
    .Z(instr_mem_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output131 (.I(net131),
    .Z(instr_mem_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output132 (.I(net132),
    .Z(instr_mem_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output133 (.I(net133),
    .Z(instr_mem_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output134 (.I(net134),
    .Z(instr_write_data[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output135 (.I(net135),
    .Z(instr_write_data[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output136 (.I(net136),
    .Z(instr_write_data[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output137 (.I(net137),
    .Z(instr_write_data[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output138 (.I(net138),
    .Z(instr_write_data[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output139 (.I(net139),
    .Z(instr_write_data[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output140 (.I(net140),
    .Z(instr_write_data[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output141 (.I(net141),
    .Z(instr_write_data[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output142 (.I(net142),
    .Z(instr_write_data[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output143 (.I(net143),
    .Z(instr_write_data[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output144 (.I(net144),
    .Z(instr_write_data[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output145 (.I(net145),
    .Z(instr_write_data[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output146 (.I(net146),
    .Z(instr_write_data[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output147 (.I(net147),
    .Z(instr_write_data[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output148 (.I(net148),
    .Z(instr_write_data[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output149 (.I(net149),
    .Z(instr_write_data[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output150 (.I(net150),
    .Z(instrw_en));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output151 (.I(net151),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output152 (.I(net152),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output153 (.I(net153),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output154 (.I(net154),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output155 (.I(net155),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output156 (.I(net156),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output157 (.I(net157),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output158 (.I(net158),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output159 (.I(net159),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output160 (.I(net160),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output161 (.I(net161),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output162 (.I(net162),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output163 (.I(net163),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output164 (.I(net164),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output165 (.I(net165),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output166 (.I(net166),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output167 (.I(net167),
    .Z(io_out[35]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output168 (.I(net168),
    .Z(la_data_out[100]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output169 (.I(net169),
    .Z(la_data_out[101]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output170 (.I(net170),
    .Z(la_data_out[102]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output171 (.I(net171),
    .Z(la_data_out[103]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output172 (.I(net172),
    .Z(la_data_out[104]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output173 (.I(net173),
    .Z(la_data_out[105]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output174 (.I(net174),
    .Z(la_data_out[106]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output175 (.I(net175),
    .Z(la_data_out[107]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output176 (.I(net176),
    .Z(la_data_out[108]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output177 (.I(net177),
    .Z(la_data_out[109]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output178 (.I(net178),
    .Z(la_data_out[110]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output179 (.I(net179),
    .Z(la_data_out[111]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output180 (.I(net180),
    .Z(la_data_out[112]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output181 (.I(net181),
    .Z(la_data_out[113]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output182 (.I(net182),
    .Z(la_data_out[114]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output183 (.I(net183),
    .Z(la_data_out[115]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output184 (.I(net184),
    .Z(la_data_out[116]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output185 (.I(net185),
    .Z(la_data_out[117]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output186 (.I(net186),
    .Z(la_data_out[118]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output187 (.I(net187),
    .Z(la_data_out[119]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output188 (.I(net188),
    .Z(la_data_out[120]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output189 (.I(net189),
    .Z(la_data_out[121]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output190 (.I(net190),
    .Z(la_data_out[122]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output191 (.I(net191),
    .Z(la_data_out[123]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output192 (.I(net192),
    .Z(la_data_out[124]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output193 (.I(net193),
    .Z(la_data_out[125]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output194 (.I(net194),
    .Z(la_data_out[126]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output195 (.I(net195),
    .Z(la_data_out[127]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output196 (.I(net196),
    .Z(la_data_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output197 (.I(net197),
    .Z(la_data_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output198 (.I(net198),
    .Z(la_data_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output199 (.I(net199),
    .Z(la_data_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output200 (.I(net200),
    .Z(la_data_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output201 (.I(net201),
    .Z(la_data_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output202 (.I(net202),
    .Z(la_data_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output203 (.I(net203),
    .Z(la_data_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output204 (.I(net204),
    .Z(la_data_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output205 (.I(net205),
    .Z(la_data_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output206 (.I(net206),
    .Z(la_data_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output207 (.I(net207),
    .Z(la_data_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output208 (.I(net208),
    .Z(la_data_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output209 (.I(net209),
    .Z(la_data_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output210 (.I(net210),
    .Z(la_data_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output211 (.I(net211),
    .Z(la_data_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output212 (.I(net212),
    .Z(la_data_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output213 (.I(net213),
    .Z(la_data_out[33]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output214 (.I(net214),
    .Z(la_data_out[34]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output215 (.I(net215),
    .Z(la_data_out[35]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output216 (.I(net216),
    .Z(la_data_out[36]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output217 (.I(net217),
    .Z(la_data_out[37]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output218 (.I(net218),
    .Z(la_data_out[38]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output219 (.I(net219),
    .Z(la_data_out[39]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output220 (.I(net220),
    .Z(la_data_out[40]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output221 (.I(net221),
    .Z(la_data_out[41]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output222 (.I(net222),
    .Z(la_data_out[42]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output223 (.I(net223),
    .Z(la_data_out[43]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output224 (.I(net224),
    .Z(la_data_out[44]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output225 (.I(net225),
    .Z(la_data_out[45]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output226 (.I(net226),
    .Z(la_data_out[46]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output227 (.I(net227),
    .Z(la_data_out[47]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output228 (.I(net228),
    .Z(la_data_out[48]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output229 (.I(net229),
    .Z(la_data_out[49]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output230 (.I(net230),
    .Z(la_data_out[50]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output231 (.I(net231),
    .Z(la_data_out[51]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output232 (.I(net232),
    .Z(la_data_out[52]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output233 (.I(net233),
    .Z(la_data_out[53]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output234 (.I(net234),
    .Z(la_data_out[54]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output235 (.I(net235),
    .Z(la_data_out[55]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output236 (.I(net236),
    .Z(la_data_out[56]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output237 (.I(net237),
    .Z(la_data_out[57]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output238 (.I(net238),
    .Z(la_data_out[58]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output239 (.I(net239),
    .Z(la_data_out[59]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output240 (.I(net240),
    .Z(la_data_out[60]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output241 (.I(net241),
    .Z(la_data_out[61]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output242 (.I(net242),
    .Z(la_data_out[62]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output243 (.I(net243),
    .Z(la_data_out[63]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output244 (.I(net244),
    .Z(la_data_out[64]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output245 (.I(net245),
    .Z(la_data_out[65]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output246 (.I(net246),
    .Z(la_data_out[66]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output247 (.I(net247),
    .Z(la_data_out[67]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output248 (.I(net248),
    .Z(la_data_out[68]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output249 (.I(net249),
    .Z(la_data_out[69]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output250 (.I(net250),
    .Z(la_data_out[70]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output251 (.I(net251),
    .Z(la_data_out[71]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output252 (.I(net252),
    .Z(la_data_out[72]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output253 (.I(net253),
    .Z(la_data_out[73]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output254 (.I(net254),
    .Z(la_data_out[74]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output255 (.I(net255),
    .Z(la_data_out[75]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output256 (.I(net256),
    .Z(la_data_out[76]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output257 (.I(net257),
    .Z(la_data_out[77]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output258 (.I(net258),
    .Z(la_data_out[78]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output259 (.I(net259),
    .Z(la_data_out[79]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output260 (.I(net260),
    .Z(la_data_out[80]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output261 (.I(net261),
    .Z(la_data_out[81]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output262 (.I(net262),
    .Z(la_data_out[82]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output263 (.I(net263),
    .Z(la_data_out[83]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output264 (.I(net264),
    .Z(la_data_out[84]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output265 (.I(net265),
    .Z(la_data_out[85]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output266 (.I(net266),
    .Z(la_data_out[86]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output267 (.I(net267),
    .Z(la_data_out[87]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output268 (.I(net268),
    .Z(la_data_out[88]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output269 (.I(net269),
    .Z(la_data_out[89]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output270 (.I(net270),
    .Z(la_data_out[90]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output271 (.I(net271),
    .Z(la_data_out[91]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output272 (.I(net272),
    .Z(la_data_out[92]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output273 (.I(net273),
    .Z(la_data_out[93]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output274 (.I(net274),
    .Z(la_data_out[94]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output275 (.I(net275),
    .Z(la_data_out[95]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output276 (.I(net276),
    .Z(la_data_out[96]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output277 (.I(net277),
    .Z(la_data_out[97]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output278 (.I(net278),
    .Z(la_data_out[98]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output279 (.I(net279),
    .Z(la_data_out[99]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output280 (.I(net280),
    .Z(reset));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output281 (.I(net281),
    .Z(start));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output282 (.I(net282),
    .Z(uP_instr[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output283 (.I(net283),
    .Z(uP_instr[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output284 (.I(net284),
    .Z(uP_instr[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output285 (.I(net285),
    .Z(uP_instr[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output286 (.I(net286),
    .Z(uP_instr[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output287 (.I(net287),
    .Z(uP_instr[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output288 (.I(net288),
    .Z(uP_instr[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output289 (.I(net289),
    .Z(uP_instr[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output290 (.I(net290),
    .Z(uP_instr[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output291 (.I(net291),
    .Z(uP_instr[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output292 (.I(net292),
    .Z(uP_instr[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output293 (.I(net293),
    .Z(uP_instr[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output294 (.I(net294),
    .Z(uP_instr[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output295 (.I(net295),
    .Z(uP_instr[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output296 (.I(net296),
    .Z(uP_instr[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output297 (.I(net297),
    .Z(uP_instr[9]));
 gf180mcu_fd_sc_mcu7t5v0__tiel io_interface_298 (.ZN(net298));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__461__A2 (.I(\Data_out0[11].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__458__A1 (.I(\Data_out0[11].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__297__I0 (.I(\Data_out0[11].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__557__B2 (.I(\Data_out0[12].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__462__A1 (.I(\Data_out0[12].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__300__I0 (.I(\Data_out0[12].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__508__B2 (.I(\Data_out0[2].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__427__A3 (.I(\Data_out0[2].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__420__A3 (.I(\Data_out0[2].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__274__I (.I(\Data_out0[2].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__512__B2 (.I(\Data_out0[3].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__393__A4 (.I(\Data_out0[3].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__390__A1 (.I(\Data_out0[3].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__256__I0 (.I(\Data_out0[3].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__511__A1 (.I(\Data_out0[3].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__427__A4 (.I(\Data_out0[3].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__424__A1 (.I(\Data_out0[3].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__279__I0 (.I(\Data_out0[3].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__523__A1 (.I(\Data_out0[5].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__398__A2 (.I(\Data_out0[5].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__397__B (.I(\Data_out0[5].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__I0 (.I(\Data_out0[5].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__526__B2 (.I(\Data_out0[5].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__433__A2 (.I(\Data_out0[5].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__432__B (.I(\Data_out0[5].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__I0 (.I(\Data_out0[5].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__531__B2 (.I(\Data_out0[6].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__402__A1 (.I(\Data_out0[6].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__401__A1 (.I(\Data_out0[6].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__I0 (.I(\Data_out0[6].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__529__I (.I(\Data_out0[6].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__442__A1 (.I(\Data_out0[6].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__534__A1 (.I(\Data_out0[7].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__405__A1 (.I(\Data_out0[7].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__266__I0 (.I(\Data_out0[7].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__535__B2 (.I(\Data_out0[7].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__442__A2 (.I(\Data_out0[7].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__441__B (.I(\Data_out0[7].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__288__I0 (.I(\Data_out0[7].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__546__B2 (.I(\Data_out0[9].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__450__A2 (.I(\Data_out0[9].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__449__B (.I(\Data_out0[9].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__I0 (.I(\Data_out0[9].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__468__A1 (.I(_023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__338__B2 (.I(_023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__331__A1 (.I(_023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__307__A1 (.I(_023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__472__I (.I(_026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__320__I (.I(_026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__I (.I(_026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__255__I (.I(_026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__473__S (.I(_027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__253__S (.I(_027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__251__S (.I(_027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__249__S (.I(_027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__556__I (.I(_030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__537__I (.I(_030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__514__I (.I(_030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__477__I (.I(_030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__485__A1 (.I(_032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__381__A1 (.I(_032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__379__A1 (.I(_032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__249__I0 (.I(_032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__534__A2 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__523__A2 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__508__A2 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__485__A2 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__511__B (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__505__B (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__497__B (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__485__B (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__567__A2 (.I(_041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__512__A2 (.I(_041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__501__A2 (.I(_041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__493__A2 (.I(_041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__557__B1 (.I(_042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__538__I (.I(_042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__507__I (.I(_042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__489__I (.I(_042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__530__A2 (.I(_043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__511__A2 (.I(_043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__497__A2 (.I(_043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__493__B1 (.I(_043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__493__B2 (.I(_044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__416__A1 (.I(_044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__413__A1 (.I(_044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__I0 (.I(_044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__567__B1 (.I(_046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__564__B1 (.I(_046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__561__B1 (.I(_046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__493__C1 (.I(_046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__502__A2 (.I(_048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__419__A1 (.I(_048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__384__A1 (.I(_048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__343__A2 (.I(_048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__497__A1 (.I(_049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__416__A2 (.I(_049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__415__A2 (.I(_049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__270__I0 (.I(_049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__501__B2 (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__389__A2 (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__381__A2 (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__251__I0 (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__502__B2 (.I(_054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__509__A2 (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__423__A1 (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__345__A2 (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__509__B1 (.I(_057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__508__A1 (.I(_058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__389__A3 (.I(_058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__386__A1 (.I(_058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__253__I0 (.I(_058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__521__A2 (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__430__A1 (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__396__A1 (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__351__A2 (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__534__B (.I(_066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__530__B (.I(_066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__523__B (.I(_066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__517__B (.I(_066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__521__B1 (.I(_067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__520__A1 (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__397__A1 (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__394__A1 (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__I0 (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__520__B2 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__432__A1 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__428__A1 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__282__I0 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__540__A2 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__535__A2 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__531__A2 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__526__A2 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__540__C1 (.I(_074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__535__C1 (.I(_074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__531__C1 (.I(_074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__526__C1 (.I(_074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__532__A2 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__440__A1 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__404__A1 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__355__A2 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__530__A1 (.I(_077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__441__A1 (.I(_077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__438__A1 (.I(_077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__286__I0 (.I(_077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__540__B2 (.I(_085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__449__A1 (.I(_085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__446__A1 (.I(_085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__291__I0 (.I(_085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__557__C1 (.I(_090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__553__C1 (.I(_090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__550__C1 (.I(_090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__546__C1 (.I(_090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__550__B2 (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__457__A1 (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__454__A1 (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__295__I0 (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__S (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__S (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__S (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__256__S (.I(_111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__299__I (.I(_116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__290__I (.I(_116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__281__I (.I(_116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__265__I (.I(_116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__271__I (.I(_120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__373__S (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__346__I (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__311__I (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__273__I (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__421__A1 (.I(_123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__278__A2 (.I(_123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__335__A1 (.I(_125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__333__A1 (.I(_125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__329__A1 (.I(_125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__277__A1 (.I(_125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__280__I (.I(_127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__362__S (.I(_138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__360__S (.I(_138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__358__S (.I(_138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__300__S (.I(_138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__327__A1 (.I(_150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__325__A1 (.I(_150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__323__A1 (.I(_150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__321__A1 (.I(_150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__363__I (.I(_173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__366__I (.I(_175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__385__I (.I(_180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__382__I (.I(_180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__377__I (.I(_180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__376__I (.I(_180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__404__B (.I(_202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__431__I (.I(_206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__422__B (.I(_206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__414__I (.I(_206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__410__I (.I(_206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__460__A1 (.I(_207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__456__A1 (.I(_207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__426__A1 (.I(_207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__413__A2 (.I(_207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__459__A2 (.I(_208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__455__A2 (.I(_208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__425__A2 (.I(_208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__412__A2 (.I(_208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__447__S (.I(_213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__439__A1 (.I(_213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__429__A1 (.I(_213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__418__B (.I(_213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__A1 (.I(_223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__453__A1 (.I(_223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__445__A1 (.I(_223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__437__A1 (.I(_223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__463__A2 (.I(_227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__452__A2 (.I(_227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__444__A2 (.I(_227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__436__A2 (.I(_227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__461__A3 (.I(_232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__451__A1 (.I(_232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__443__I (.I(_232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__457__A2 (.I(_233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__449__A2 (.I(_233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__446__A2 (.I(_233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__445__A3 (.I(_233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(data_read_data[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(data_read_data[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(data_read_data[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(data_read_data[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(data_read_data[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(data_read_data[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(data_read_data[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(data_read_data[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(data_read_data[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(data_read_data[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(data_read_data[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(data_read_data[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(data_read_data[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(data_read_data[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(data_read_data[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(data_read_data[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(hlt));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(instr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(instr[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(instr[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(instr[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(instr[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(instr[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(instr[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(instr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(instr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(instr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(instr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(instr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(instr[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(instr[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(instr[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(instr[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(io_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(io_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(io_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(io_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(io_in[32]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(io_in[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(io_in[34]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(io_in[36]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(io_in[37]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(uP_data_mem_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(uP_data_mem_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(uP_data_mem_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(uP_data_mem_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(uP_data_mem_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(uP_data_mem_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(uP_data_mem_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(uP_data_mem_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(uP_dataw_en));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(uP_instr_mem_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(uP_instr_mem_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(uP_instr_mem_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(uP_instr_mem_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(uP_instr_mem_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(uP_instr_mem_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(uP_instr_mem_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(uP_instr_mem_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(uP_instr_mem_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input73_I (.I(uP_instr_mem_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input74_I (.I(uP_instr_mem_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input75_I (.I(uP_instr_mem_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input76_I (.I(uP_instr_mem_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input77_I (.I(uP_write_data[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input78_I (.I(uP_write_data[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input79_I (.I(uP_write_data[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input80_I (.I(uP_write_data[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input81_I (.I(uP_write_data[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input82_I (.I(uP_write_data[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input83_I (.I(uP_write_data[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input84_I (.I(uP_write_data[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input85_I (.I(uP_write_data[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input86_I (.I(uP_write_data[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input87_I (.I(uP_write_data[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input88_I (.I(uP_write_data[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input89_I (.I(uP_write_data[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input90_I (.I(uP_write_data[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input91_I (.I(uP_write_data[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input92_I (.I(uP_write_data[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input93_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input94_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__715__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__493__C2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__725__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__550__C2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__726__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__553__C2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__727__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__557__C2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__728__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__561__B2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__729__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__564__B2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__730__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__567__B2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__716__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__501__C2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__717__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__508__C2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__718__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__512__C2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__719__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__520__C2 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__720__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__526__C2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__721__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__531__C2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__722__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__535__C2 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__723__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__540__C2 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__724__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__546__C2 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__685__I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__493__A1 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__303__A2 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__550__A1 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__325__A2 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__553__A1 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__327__A2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__557__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__329__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__561__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__331__A2 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__564__A1 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__333__A2 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__567__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__335__A2 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__501__A1 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__305__A2 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__505__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__307__A2 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__512__A1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__309__A2 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__517__A1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__312__A2 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__526__A1 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__314__A2 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__531__A1 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__316__A2 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__535__A1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__318__A2 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__540__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__321__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__546__A1 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__323__A2 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__758__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__669__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__475__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__412__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__378__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__768__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__679__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__551__A2 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__455__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__362__I0 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__769__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__680__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__554__A2 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__459__A1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__365__I0 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__770__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__681__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__559__A2 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__463__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__367__I0 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__771__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__682__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__562__A2 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__369__I0 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__772__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__683__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__565__A2 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__371__I0 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__773__I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__684__I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__568__A2 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__373__I0 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__759__I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__670__I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__495__I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__760__I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__671__I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__503__I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__387__A1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__755__I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__483__I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__476__I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__468__A2 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__756__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__480__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__466__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__757__I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__479__I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__465__I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__783__I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__774__I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__470__I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__467__I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__779__I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__473__I0 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__761__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__672__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__510__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__425__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__391__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__762__I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__673__I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__515__I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__763__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__674__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__522__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__436__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__399__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__764__I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__675__I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__528__I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__765__I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__676__I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__533__I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__444__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__406__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__766__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__677__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__542__A2 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__447__I1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__358__I0 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__767__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__678__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__547__A2 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__452__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__360__I0 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__249__I1 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__251__I1 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__253__I1 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__256__I1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__I1 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__I1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__I1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__266__I1 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__777__I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__337__I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__I1 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__295__I1 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__297__I1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__300__I1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__270__I1 (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__277__A2 (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__279__I1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__282__I1 (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__I1 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__286__I1 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__288__I1 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__291__I1 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__I1 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__780__I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__473__I1 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__782__I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__778__I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__590__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__589__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__588__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__587__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__586__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__585__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__584__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__583__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__582__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__581__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__580__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__579__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__578__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__577__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__576__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__575__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__574__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__573__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__572__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__571__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__570__RN (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output95_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__781__I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__590__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__589__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__588__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__587__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__586__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__585__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__584__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__583__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__582__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__581__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__580__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__579__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__578__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__577__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__576__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__575__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__574__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__573__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__572__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__571__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__570__CLK (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output96_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__731__I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output97_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__732__I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output98_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__733__I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output99_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__734__I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output100_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__735__I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output101_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__736__I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output102_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__737__I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output103_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__738__I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output104_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__699__I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output105_I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__709__I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output106_I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__710__I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output107_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__711__I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output108_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__712__I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output109_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__713__I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output110_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__714__I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output111_I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__700__I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output112_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__701__I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output113_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__702__I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output114_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__703__I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output115_I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__704__I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output116_I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__705__I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output117_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__706__I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output118_I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__707__I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output119_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__708__I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output120_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__776__I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output121_I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__686__I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output122_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__696__I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output123_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__697__I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output124_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__698__I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output125_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__687__I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output126_I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__688__I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output127_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__689__I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output128_I (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__690__I (.I(net128));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output129_I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__691__I (.I(net129));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output130_I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__692__I (.I(net130));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output131_I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__693__I (.I(net131));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output132_I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__694__I (.I(net132));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output133_I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__695__I (.I(net133));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output135_I (.I(net135));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output136_I (.I(net136));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output137_I (.I(net137));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output138_I (.I(net138));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output139_I (.I(net139));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output140_I (.I(net140));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output143_I (.I(net143));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output145_I (.I(net145));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output148_I (.I(net148));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output149_I (.I(net149));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output150_I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__775__I (.I(net150));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output151_I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__739__I (.I(net151));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output152_I (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__740__I (.I(net152));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output153_I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__741__I (.I(net153));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output154_I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__742__I (.I(net154));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output155_I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__743__I (.I(net155));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output156_I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__744__I (.I(net156));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output157_I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__745__I (.I(net157));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output158_I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__746__I (.I(net158));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output159_I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__747__I (.I(net159));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output160_I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__748__I (.I(net160));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output161_I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__749__I (.I(net161));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output162_I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__750__I (.I(net162));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output163_I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__751__I (.I(net163));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output164_I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__752__I (.I(net164));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output165_I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__753__I (.I(net165));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output166_I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__754__I (.I(net166));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output168_I (.I(net168));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output169_I (.I(net169));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output170_I (.I(net170));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output171_I (.I(net171));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output174_I (.I(net174));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output175_I (.I(net175));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output176_I (.I(net176));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output179_I (.I(net179));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output180_I (.I(net180));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output181_I (.I(net181));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output182_I (.I(net182));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output183_I (.I(net183));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output184_I (.I(net184));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output185_I (.I(net185));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output186_I (.I(net186));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output187_I (.I(net187));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output189_I (.I(net189));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output190_I (.I(net190));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output191_I (.I(net191));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output193_I (.I(net193));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output196_I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__784__I (.I(net196));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output197_I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__785__I (.I(net197));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output198_I (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__786__I (.I(net198));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output199_I (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__787__I (.I(net199));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output200_I (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__788__I (.I(net200));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output201_I (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__789__I (.I(net201));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output202_I (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__790__I (.I(net202));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output203_I (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__791__I (.I(net203));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output204_I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__792__I (.I(net204));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output205_I (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__793__I (.I(net205));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output206_I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__794__I (.I(net206));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output207_I (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__795__I (.I(net207));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output208_I (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__796__I (.I(net208));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output209_I (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__797__I (.I(net209));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output210_I (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__798__I (.I(net210));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output211_I (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__799__I (.I(net211));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output212_I (.I(net212));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output213_I (.I(net213));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output214_I (.I(net214));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output215_I (.I(net215));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output216_I (.I(net216));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output217_I (.I(net217));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output218_I (.I(net218));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output219_I (.I(net219));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output220_I (.I(net220));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output221_I (.I(net221));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output222_I (.I(net222));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output223_I (.I(net223));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output224_I (.I(net224));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output225_I (.I(net225));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output226_I (.I(net226));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output227_I (.I(net227));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output228_I (.I(net228));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output229_I (.I(net229));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output230_I (.I(net230));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output231_I (.I(net231));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output232_I (.I(net232));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output233_I (.I(net233));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output234_I (.I(net234));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output235_I (.I(net235));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output236_I (.I(net236));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output237_I (.I(net237));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output238_I (.I(net238));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output239_I (.I(net239));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output240_I (.I(net240));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output241_I (.I(net241));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output242_I (.I(net242));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output243_I (.I(net243));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output244_I (.I(net244));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output245_I (.I(net245));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output246_I (.I(net246));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output247_I (.I(net247));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output248_I (.I(net248));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output249_I (.I(net249));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output250_I (.I(net250));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output251_I (.I(net251));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output252_I (.I(net252));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output253_I (.I(net253));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output254_I (.I(net254));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output255_I (.I(net255));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output256_I (.I(net256));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output257_I (.I(net257));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output258_I (.I(net258));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output259_I (.I(net259));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output260_I (.I(net260));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output261_I (.I(net261));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output262_I (.I(net262));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output263_I (.I(net263));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output264_I (.I(net264));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output265_I (.I(net265));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output266_I (.I(net266));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output267_I (.I(net267));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output268_I (.I(net268));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output269_I (.I(net269));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output270_I (.I(net270));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output271_I (.I(net271));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output272_I (.I(net272));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output273_I (.I(net273));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output274_I (.I(net274));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output275_I (.I(net275));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output276_I (.I(net276));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output277_I (.I(net277));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output278_I (.I(net278));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output279_I (.I(net279));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output280_I (.I(net280));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output281_I (.I(net281));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output282_I (.I(net282));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output289_I (.I(net289));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output290_I (.I(net290));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output292_I (.I(net292));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1044 ();
 assign io_oeb[0] = net355;
 assign io_oeb[10] = net365;
 assign io_oeb[11] = net366;
 assign io_oeb[12] = net367;
 assign io_oeb[13] = net368;
 assign io_oeb[14] = net369;
 assign io_oeb[15] = net370;
 assign io_oeb[16] = net298;
 assign io_oeb[17] = net299;
 assign io_oeb[18] = net300;
 assign io_oeb[19] = net301;
 assign io_oeb[1] = net356;
 assign io_oeb[20] = net302;
 assign io_oeb[21] = net303;
 assign io_oeb[22] = net304;
 assign io_oeb[23] = net305;
 assign io_oeb[24] = net306;
 assign io_oeb[25] = net307;
 assign io_oeb[26] = net308;
 assign io_oeb[27] = net309;
 assign io_oeb[28] = net310;
 assign io_oeb[29] = net311;
 assign io_oeb[2] = net357;
 assign io_oeb[30] = net312;
 assign io_oeb[31] = net313;
 assign io_oeb[32] = net371;
 assign io_oeb[33] = net372;
 assign io_oeb[34] = net373;
 assign io_oeb[35] = net314;
 assign io_oeb[36] = net374;
 assign io_oeb[37] = net375;
 assign io_oeb[3] = net358;
 assign io_oeb[4] = net359;
 assign io_oeb[5] = net360;
 assign io_oeb[6] = net361;
 assign io_oeb[7] = net362;
 assign io_oeb[8] = net363;
 assign io_oeb[9] = net364;
 assign io_out[0] = net315;
 assign io_out[10] = net325;
 assign io_out[11] = net326;
 assign io_out[12] = net327;
 assign io_out[13] = net328;
 assign io_out[14] = net329;
 assign io_out[15] = net330;
 assign io_out[1] = net316;
 assign io_out[2] = net317;
 assign io_out[32] = net331;
 assign io_out[33] = net332;
 assign io_out[34] = net333;
 assign io_out[36] = net334;
 assign io_out[37] = net335;
 assign io_out[3] = net318;
 assign io_out[4] = net319;
 assign io_out[5] = net320;
 assign io_out[6] = net321;
 assign io_out[7] = net322;
 assign io_out[8] = net323;
 assign io_out[9] = net324;
 assign irq[0] = net336;
 assign irq[1] = net337;
 assign irq[2] = net338;
 assign la_data_out[0] = net339;
 assign la_data_out[10] = net349;
 assign la_data_out[11] = net350;
 assign la_data_out[12] = net351;
 assign la_data_out[13] = net352;
 assign la_data_out[14] = net353;
 assign la_data_out[15] = net354;
 assign la_data_out[1] = net340;
 assign la_data_out[2] = net341;
 assign la_data_out[3] = net342;
 assign la_data_out[4] = net343;
 assign la_data_out[5] = net344;
 assign la_data_out[6] = net345;
 assign la_data_out[7] = net346;
 assign la_data_out[8] = net347;
 assign la_data_out[9] = net348;
endmodule

