VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO processor
  CLASS BLOCK ;
  FOREIGN processor ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 1000.000 ;
  PIN Dataw_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 943.040 996.000 943.600 1000.000 ;
    END
  END Dataw_en
  PIN Serial_input
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 969.920 996.000 970.480 1000.000 ;
    END
  END Serial_input
  PIN Serial_output
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 983.360 996.000 983.920 1000.000 ;
    END
  END Serial_output
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 166.320 0.000 166.880 4.000 ;
    END
  END clk
  PIN data_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 405.440 996.000 406.000 1000.000 ;
    END
  END data_mem_addr[0]
  PIN data_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 418.880 996.000 419.440 1000.000 ;
    END
  END data_mem_addr[1]
  PIN data_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 432.320 996.000 432.880 1000.000 ;
    END
  END data_mem_addr[2]
  PIN data_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 445.760 996.000 446.320 1000.000 ;
    END
  END data_mem_addr[3]
  PIN data_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 459.200 996.000 459.760 1000.000 ;
    END
  END data_mem_addr[4]
  PIN data_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 472.640 996.000 473.200 1000.000 ;
    END
  END data_mem_addr[5]
  PIN data_mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 486.080 996.000 486.640 1000.000 ;
    END
  END data_mem_addr[6]
  PIN data_mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 499.520 996.000 500.080 1000.000 ;
    END
  END data_mem_addr[7]
  PIN hlt
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 956.480 996.000 957.040 1000.000 ;
    END
  END hlt
  PIN instr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 15.680 996.000 16.240 1000.000 ;
    END
  END instr[0]
  PIN instr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 284.480 996.000 285.040 1000.000 ;
    END
  END instr[10]
  PIN instr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 311.360 996.000 311.920 1000.000 ;
    END
  END instr[11]
  PIN instr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 338.240 996.000 338.800 1000.000 ;
    END
  END instr[12]
  PIN instr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 365.120 996.000 365.680 1000.000 ;
    END
  END instr[13]
  PIN instr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 378.560 996.000 379.120 1000.000 ;
    END
  END instr[14]
  PIN instr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 392.000 996.000 392.560 1000.000 ;
    END
  END instr[15]
  PIN instr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 42.560 996.000 43.120 1000.000 ;
    END
  END instr[1]
  PIN instr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 996.000 70.000 1000.000 ;
    END
  END instr[2]
  PIN instr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 996.000 96.880 1000.000 ;
    END
  END instr[3]
  PIN instr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 996.000 123.760 1000.000 ;
    END
  END instr[4]
  PIN instr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 150.080 996.000 150.640 1000.000 ;
    END
  END instr[5]
  PIN instr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 176.960 996.000 177.520 1000.000 ;
    END
  END instr[6]
  PIN instr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 203.840 996.000 204.400 1000.000 ;
    END
  END instr[7]
  PIN instr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 230.720 996.000 231.280 1000.000 ;
    END
  END instr[8]
  PIN instr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 257.600 996.000 258.160 1000.000 ;
    END
  END instr[9]
  PIN instr_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.120 996.000 29.680 1000.000 ;
    END
  END instr_mem_addr[0]
  PIN instr_mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 297.920 996.000 298.480 1000.000 ;
    END
  END instr_mem_addr[10]
  PIN instr_mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 324.800 996.000 325.360 1000.000 ;
    END
  END instr_mem_addr[11]
  PIN instr_mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 351.680 996.000 352.240 1000.000 ;
    END
  END instr_mem_addr[12]
  PIN instr_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 56.000 996.000 56.560 1000.000 ;
    END
  END instr_mem_addr[1]
  PIN instr_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 82.880 996.000 83.440 1000.000 ;
    END
  END instr_mem_addr[2]
  PIN instr_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 109.760 996.000 110.320 1000.000 ;
    END
  END instr_mem_addr[3]
  PIN instr_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 136.640 996.000 137.200 1000.000 ;
    END
  END instr_mem_addr[4]
  PIN instr_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 163.520 996.000 164.080 1000.000 ;
    END
  END instr_mem_addr[5]
  PIN instr_mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 190.400 996.000 190.960 1000.000 ;
    END
  END instr_mem_addr[6]
  PIN instr_mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 217.280 996.000 217.840 1000.000 ;
    END
  END instr_mem_addr[7]
  PIN instr_mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 244.160 996.000 244.720 1000.000 ;
    END
  END instr_mem_addr[8]
  PIN instr_mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 271.040 996.000 271.600 1000.000 ;
    END
  END instr_mem_addr[9]
  PIN read_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 512.960 996.000 513.520 1000.000 ;
    END
  END read_data[0]
  PIN read_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 647.360 996.000 647.920 1000.000 ;
    END
  END read_data[10]
  PIN read_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 660.800 996.000 661.360 1000.000 ;
    END
  END read_data[11]
  PIN read_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 674.240 996.000 674.800 1000.000 ;
    END
  END read_data[12]
  PIN read_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 687.680 996.000 688.240 1000.000 ;
    END
  END read_data[13]
  PIN read_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 701.120 996.000 701.680 1000.000 ;
    END
  END read_data[14]
  PIN read_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 714.560 996.000 715.120 1000.000 ;
    END
  END read_data[15]
  PIN read_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 526.400 996.000 526.960 1000.000 ;
    END
  END read_data[1]
  PIN read_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 539.840 996.000 540.400 1000.000 ;
    END
  END read_data[2]
  PIN read_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 553.280 996.000 553.840 1000.000 ;
    END
  END read_data[3]
  PIN read_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 566.720 996.000 567.280 1000.000 ;
    END
  END read_data[4]
  PIN read_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 580.160 996.000 580.720 1000.000 ;
    END
  END read_data[5]
  PIN read_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 593.600 996.000 594.160 1000.000 ;
    END
  END read_data[6]
  PIN read_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 607.040 996.000 607.600 1000.000 ;
    END
  END read_data[7]
  PIN read_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 620.480 996.000 621.040 1000.000 ;
    END
  END read_data[8]
  PIN read_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 633.920 996.000 634.480 1000.000 ;
    END
  END read_data[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 499.520 0.000 500.080 4.000 ;
    END
  END reset
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 832.720 0.000 833.280 4.000 ;
    END
  END start
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 984.220 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 984.220 ;
    END
  END vss
  PIN write_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 728.000 996.000 728.560 1000.000 ;
    END
  END write_data[0]
  PIN write_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 862.400 996.000 862.960 1000.000 ;
    END
  END write_data[10]
  PIN write_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 875.840 996.000 876.400 1000.000 ;
    END
  END write_data[11]
  PIN write_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 889.280 996.000 889.840 1000.000 ;
    END
  END write_data[12]
  PIN write_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 902.720 996.000 903.280 1000.000 ;
    END
  END write_data[13]
  PIN write_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 916.160 996.000 916.720 1000.000 ;
    END
  END write_data[14]
  PIN write_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 929.600 996.000 930.160 1000.000 ;
    END
  END write_data[15]
  PIN write_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 741.440 996.000 742.000 1000.000 ;
    END
  END write_data[1]
  PIN write_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 754.880 996.000 755.440 1000.000 ;
    END
  END write_data[2]
  PIN write_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 768.320 996.000 768.880 1000.000 ;
    END
  END write_data[3]
  PIN write_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 781.760 996.000 782.320 1000.000 ;
    END
  END write_data[4]
  PIN write_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 795.200 996.000 795.760 1000.000 ;
    END
  END write_data[5]
  PIN write_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 808.640 996.000 809.200 1000.000 ;
    END
  END write_data[6]
  PIN write_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 822.080 996.000 822.640 1000.000 ;
    END
  END write_data[7]
  PIN write_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 835.520 996.000 836.080 1000.000 ;
    END
  END write_data[8]
  PIN write_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 848.960 996.000 849.520 1000.000 ;
    END
  END write_data[9]
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 992.880 984.220 ;
      LAYER Metal2 ;
        RECT 14.700 995.700 15.380 996.660 ;
        RECT 16.540 995.700 28.820 996.660 ;
        RECT 29.980 995.700 42.260 996.660 ;
        RECT 43.420 995.700 55.700 996.660 ;
        RECT 56.860 995.700 69.140 996.660 ;
        RECT 70.300 995.700 82.580 996.660 ;
        RECT 83.740 995.700 96.020 996.660 ;
        RECT 97.180 995.700 109.460 996.660 ;
        RECT 110.620 995.700 122.900 996.660 ;
        RECT 124.060 995.700 136.340 996.660 ;
        RECT 137.500 995.700 149.780 996.660 ;
        RECT 150.940 995.700 163.220 996.660 ;
        RECT 164.380 995.700 176.660 996.660 ;
        RECT 177.820 995.700 190.100 996.660 ;
        RECT 191.260 995.700 203.540 996.660 ;
        RECT 204.700 995.700 216.980 996.660 ;
        RECT 218.140 995.700 230.420 996.660 ;
        RECT 231.580 995.700 243.860 996.660 ;
        RECT 245.020 995.700 257.300 996.660 ;
        RECT 258.460 995.700 270.740 996.660 ;
        RECT 271.900 995.700 284.180 996.660 ;
        RECT 285.340 995.700 297.620 996.660 ;
        RECT 298.780 995.700 311.060 996.660 ;
        RECT 312.220 995.700 324.500 996.660 ;
        RECT 325.660 995.700 337.940 996.660 ;
        RECT 339.100 995.700 351.380 996.660 ;
        RECT 352.540 995.700 364.820 996.660 ;
        RECT 365.980 995.700 378.260 996.660 ;
        RECT 379.420 995.700 391.700 996.660 ;
        RECT 392.860 995.700 405.140 996.660 ;
        RECT 406.300 995.700 418.580 996.660 ;
        RECT 419.740 995.700 432.020 996.660 ;
        RECT 433.180 995.700 445.460 996.660 ;
        RECT 446.620 995.700 458.900 996.660 ;
        RECT 460.060 995.700 472.340 996.660 ;
        RECT 473.500 995.700 485.780 996.660 ;
        RECT 486.940 995.700 499.220 996.660 ;
        RECT 500.380 995.700 512.660 996.660 ;
        RECT 513.820 995.700 526.100 996.660 ;
        RECT 527.260 995.700 539.540 996.660 ;
        RECT 540.700 995.700 552.980 996.660 ;
        RECT 554.140 995.700 566.420 996.660 ;
        RECT 567.580 995.700 579.860 996.660 ;
        RECT 581.020 995.700 593.300 996.660 ;
        RECT 594.460 995.700 606.740 996.660 ;
        RECT 607.900 995.700 620.180 996.660 ;
        RECT 621.340 995.700 633.620 996.660 ;
        RECT 634.780 995.700 647.060 996.660 ;
        RECT 648.220 995.700 660.500 996.660 ;
        RECT 661.660 995.700 673.940 996.660 ;
        RECT 675.100 995.700 687.380 996.660 ;
        RECT 688.540 995.700 700.820 996.660 ;
        RECT 701.980 995.700 714.260 996.660 ;
        RECT 715.420 995.700 727.700 996.660 ;
        RECT 728.860 995.700 741.140 996.660 ;
        RECT 742.300 995.700 754.580 996.660 ;
        RECT 755.740 995.700 768.020 996.660 ;
        RECT 769.180 995.700 781.460 996.660 ;
        RECT 782.620 995.700 794.900 996.660 ;
        RECT 796.060 995.700 808.340 996.660 ;
        RECT 809.500 995.700 821.780 996.660 ;
        RECT 822.940 995.700 835.220 996.660 ;
        RECT 836.380 995.700 848.660 996.660 ;
        RECT 849.820 995.700 862.100 996.660 ;
        RECT 863.260 995.700 875.540 996.660 ;
        RECT 876.700 995.700 888.980 996.660 ;
        RECT 890.140 995.700 902.420 996.660 ;
        RECT 903.580 995.700 915.860 996.660 ;
        RECT 917.020 995.700 929.300 996.660 ;
        RECT 930.460 995.700 942.740 996.660 ;
        RECT 943.900 995.700 956.180 996.660 ;
        RECT 957.340 995.700 969.620 996.660 ;
        RECT 970.780 995.700 983.060 996.660 ;
        RECT 14.700 4.300 983.780 995.700 ;
        RECT 14.700 4.000 166.020 4.300 ;
        RECT 167.180 4.000 499.220 4.300 ;
        RECT 500.380 4.000 832.420 4.300 ;
        RECT 833.580 4.000 983.780 4.300 ;
      LAYER Metal3 ;
        RECT 18.570 15.540 979.350 985.460 ;
      LAYER Metal4 ;
        RECT 251.580 545.530 252.340 973.190 ;
        RECT 254.540 545.530 329.140 973.190 ;
        RECT 331.340 545.530 405.940 973.190 ;
        RECT 408.140 545.530 482.740 973.190 ;
        RECT 484.940 545.530 559.540 973.190 ;
        RECT 561.740 545.530 636.340 973.190 ;
        RECT 638.540 545.530 713.140 973.190 ;
        RECT 715.340 545.530 776.580 973.190 ;
  END
END processor
END LIBRARY

