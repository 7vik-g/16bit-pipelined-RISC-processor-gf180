magic
tech gf180mcuC
magscale 1 5
timestamp 1670663505
<< obsm1 >>
rect 672 1415 179312 98489
<< metal2 >>
rect 6776 99600 6832 100000
rect 7392 99600 7448 100000
rect 8008 99600 8064 100000
rect 8624 99600 8680 100000
rect 9240 99600 9296 100000
rect 9856 99600 9912 100000
rect 10472 99600 10528 100000
rect 11088 99600 11144 100000
rect 11704 99600 11760 100000
rect 12320 99600 12376 100000
rect 12936 99600 12992 100000
rect 13552 99600 13608 100000
rect 14168 99600 14224 100000
rect 14784 99600 14840 100000
rect 15400 99600 15456 100000
rect 16016 99600 16072 100000
rect 16632 99600 16688 100000
rect 17248 99600 17304 100000
rect 17864 99600 17920 100000
rect 18480 99600 18536 100000
rect 19096 99600 19152 100000
rect 19712 99600 19768 100000
rect 20328 99600 20384 100000
rect 20944 99600 21000 100000
rect 21560 99600 21616 100000
rect 22176 99600 22232 100000
rect 22792 99600 22848 100000
rect 23408 99600 23464 100000
rect 24024 99600 24080 100000
rect 24640 99600 24696 100000
rect 25256 99600 25312 100000
rect 25872 99600 25928 100000
rect 26488 99600 26544 100000
rect 27104 99600 27160 100000
rect 27720 99600 27776 100000
rect 28336 99600 28392 100000
rect 28952 99600 29008 100000
rect 29568 99600 29624 100000
rect 30184 99600 30240 100000
rect 30800 99600 30856 100000
rect 31416 99600 31472 100000
rect 32032 99600 32088 100000
rect 32648 99600 32704 100000
rect 33264 99600 33320 100000
rect 33880 99600 33936 100000
rect 34496 99600 34552 100000
rect 35112 99600 35168 100000
rect 35728 99600 35784 100000
rect 36344 99600 36400 100000
rect 36960 99600 37016 100000
rect 37576 99600 37632 100000
rect 38192 99600 38248 100000
rect 38808 99600 38864 100000
rect 39424 99600 39480 100000
rect 40040 99600 40096 100000
rect 40656 99600 40712 100000
rect 41272 99600 41328 100000
rect 41888 99600 41944 100000
rect 42504 99600 42560 100000
rect 43120 99600 43176 100000
rect 43736 99600 43792 100000
rect 44352 99600 44408 100000
rect 44968 99600 45024 100000
rect 45584 99600 45640 100000
rect 46200 99600 46256 100000
rect 46816 99600 46872 100000
rect 47432 99600 47488 100000
rect 48048 99600 48104 100000
rect 48664 99600 48720 100000
rect 49280 99600 49336 100000
rect 49896 99600 49952 100000
rect 50512 99600 50568 100000
rect 51128 99600 51184 100000
rect 51744 99600 51800 100000
rect 52360 99600 52416 100000
rect 52976 99600 53032 100000
rect 53592 99600 53648 100000
rect 54208 99600 54264 100000
rect 54824 99600 54880 100000
rect 55440 99600 55496 100000
rect 56056 99600 56112 100000
rect 56672 99600 56728 100000
rect 57288 99600 57344 100000
rect 57904 99600 57960 100000
rect 58520 99600 58576 100000
rect 59136 99600 59192 100000
rect 59752 99600 59808 100000
rect 60368 99600 60424 100000
rect 60984 99600 61040 100000
rect 61600 99600 61656 100000
rect 62216 99600 62272 100000
rect 62832 99600 62888 100000
rect 63448 99600 63504 100000
rect 64064 99600 64120 100000
rect 64680 99600 64736 100000
rect 65296 99600 65352 100000
rect 65912 99600 65968 100000
rect 66528 99600 66584 100000
rect 67144 99600 67200 100000
rect 67760 99600 67816 100000
rect 68376 99600 68432 100000
rect 68992 99600 69048 100000
rect 69608 99600 69664 100000
rect 70224 99600 70280 100000
rect 70840 99600 70896 100000
rect 71456 99600 71512 100000
rect 72072 99600 72128 100000
rect 72688 99600 72744 100000
rect 73304 99600 73360 100000
rect 73920 99600 73976 100000
rect 74536 99600 74592 100000
rect 75152 99600 75208 100000
rect 75768 99600 75824 100000
rect 76384 99600 76440 100000
rect 77000 99600 77056 100000
rect 77616 99600 77672 100000
rect 78232 99600 78288 100000
rect 78848 99600 78904 100000
rect 79464 99600 79520 100000
rect 80080 99600 80136 100000
rect 80696 99600 80752 100000
rect 81312 99600 81368 100000
rect 81928 99600 81984 100000
rect 82544 99600 82600 100000
rect 83160 99600 83216 100000
rect 83776 99600 83832 100000
rect 84392 99600 84448 100000
rect 85008 99600 85064 100000
rect 85624 99600 85680 100000
rect 86240 99600 86296 100000
rect 86856 99600 86912 100000
rect 87472 99600 87528 100000
rect 88088 99600 88144 100000
rect 88704 99600 88760 100000
rect 89320 99600 89376 100000
rect 89936 99600 89992 100000
rect 90552 99600 90608 100000
rect 91168 99600 91224 100000
rect 91784 99600 91840 100000
rect 92400 99600 92456 100000
rect 93016 99600 93072 100000
rect 93632 99600 93688 100000
rect 94248 99600 94304 100000
rect 94864 99600 94920 100000
rect 95480 99600 95536 100000
rect 96096 99600 96152 100000
rect 96712 99600 96768 100000
rect 97328 99600 97384 100000
rect 97944 99600 98000 100000
rect 98560 99600 98616 100000
rect 99176 99600 99232 100000
rect 99792 99600 99848 100000
rect 100408 99600 100464 100000
rect 101024 99600 101080 100000
rect 101640 99600 101696 100000
rect 102256 99600 102312 100000
rect 102872 99600 102928 100000
rect 103488 99600 103544 100000
rect 104104 99600 104160 100000
rect 104720 99600 104776 100000
rect 105336 99600 105392 100000
rect 105952 99600 106008 100000
rect 106568 99600 106624 100000
rect 107184 99600 107240 100000
rect 107800 99600 107856 100000
rect 108416 99600 108472 100000
rect 109032 99600 109088 100000
rect 109648 99600 109704 100000
rect 110264 99600 110320 100000
rect 110880 99600 110936 100000
rect 111496 99600 111552 100000
rect 112112 99600 112168 100000
rect 112728 99600 112784 100000
rect 113344 99600 113400 100000
rect 113960 99600 114016 100000
rect 114576 99600 114632 100000
rect 115192 99600 115248 100000
rect 115808 99600 115864 100000
rect 116424 99600 116480 100000
rect 117040 99600 117096 100000
rect 117656 99600 117712 100000
rect 118272 99600 118328 100000
rect 118888 99600 118944 100000
rect 119504 99600 119560 100000
rect 120120 99600 120176 100000
rect 120736 99600 120792 100000
rect 121352 99600 121408 100000
rect 121968 99600 122024 100000
rect 122584 99600 122640 100000
rect 123200 99600 123256 100000
rect 123816 99600 123872 100000
rect 124432 99600 124488 100000
rect 125048 99600 125104 100000
rect 125664 99600 125720 100000
rect 126280 99600 126336 100000
rect 126896 99600 126952 100000
rect 127512 99600 127568 100000
rect 128128 99600 128184 100000
rect 128744 99600 128800 100000
rect 129360 99600 129416 100000
rect 129976 99600 130032 100000
rect 130592 99600 130648 100000
rect 131208 99600 131264 100000
rect 131824 99600 131880 100000
rect 132440 99600 132496 100000
rect 133056 99600 133112 100000
rect 133672 99600 133728 100000
rect 134288 99600 134344 100000
rect 134904 99600 134960 100000
rect 135520 99600 135576 100000
rect 136136 99600 136192 100000
rect 136752 99600 136808 100000
rect 137368 99600 137424 100000
rect 137984 99600 138040 100000
rect 138600 99600 138656 100000
rect 139216 99600 139272 100000
rect 139832 99600 139888 100000
rect 140448 99600 140504 100000
rect 141064 99600 141120 100000
rect 141680 99600 141736 100000
rect 142296 99600 142352 100000
rect 142912 99600 142968 100000
rect 143528 99600 143584 100000
rect 144144 99600 144200 100000
rect 144760 99600 144816 100000
rect 145376 99600 145432 100000
rect 145992 99600 146048 100000
rect 146608 99600 146664 100000
rect 147224 99600 147280 100000
rect 147840 99600 147896 100000
rect 148456 99600 148512 100000
rect 149072 99600 149128 100000
rect 149688 99600 149744 100000
rect 150304 99600 150360 100000
rect 150920 99600 150976 100000
rect 151536 99600 151592 100000
rect 152152 99600 152208 100000
rect 152768 99600 152824 100000
rect 153384 99600 153440 100000
rect 154000 99600 154056 100000
rect 154616 99600 154672 100000
rect 155232 99600 155288 100000
rect 155848 99600 155904 100000
rect 156464 99600 156520 100000
rect 157080 99600 157136 100000
rect 157696 99600 157752 100000
rect 158312 99600 158368 100000
rect 158928 99600 158984 100000
rect 159544 99600 159600 100000
rect 160160 99600 160216 100000
rect 160776 99600 160832 100000
rect 161392 99600 161448 100000
rect 162008 99600 162064 100000
rect 162624 99600 162680 100000
rect 163240 99600 163296 100000
rect 163856 99600 163912 100000
rect 164472 99600 164528 100000
rect 165088 99600 165144 100000
rect 165704 99600 165760 100000
rect 166320 99600 166376 100000
rect 166936 99600 166992 100000
rect 167552 99600 167608 100000
rect 168168 99600 168224 100000
rect 168784 99600 168840 100000
rect 169400 99600 169456 100000
rect 170016 99600 170072 100000
rect 170632 99600 170688 100000
rect 171248 99600 171304 100000
rect 171864 99600 171920 100000
rect 172480 99600 172536 100000
rect 173096 99600 173152 100000
rect 1904 0 1960 400
rect 2240 0 2296 400
rect 2576 0 2632 400
rect 2912 0 2968 400
rect 3248 0 3304 400
rect 3584 0 3640 400
rect 3920 0 3976 400
rect 4256 0 4312 400
rect 4592 0 4648 400
rect 4928 0 4984 400
rect 5264 0 5320 400
rect 5600 0 5656 400
rect 5936 0 5992 400
rect 6272 0 6328 400
rect 6608 0 6664 400
rect 6944 0 7000 400
rect 7280 0 7336 400
rect 7616 0 7672 400
rect 7952 0 8008 400
rect 8288 0 8344 400
rect 8624 0 8680 400
rect 8960 0 9016 400
rect 9296 0 9352 400
rect 9632 0 9688 400
rect 9968 0 10024 400
rect 10304 0 10360 400
rect 10640 0 10696 400
rect 10976 0 11032 400
rect 11312 0 11368 400
rect 11648 0 11704 400
rect 11984 0 12040 400
rect 12320 0 12376 400
rect 12656 0 12712 400
rect 12992 0 13048 400
rect 13328 0 13384 400
rect 13664 0 13720 400
rect 14000 0 14056 400
rect 14336 0 14392 400
rect 14672 0 14728 400
rect 15008 0 15064 400
rect 15344 0 15400 400
rect 15680 0 15736 400
rect 16016 0 16072 400
rect 16352 0 16408 400
rect 16688 0 16744 400
rect 17024 0 17080 400
rect 17360 0 17416 400
rect 17696 0 17752 400
rect 18032 0 18088 400
rect 18368 0 18424 400
rect 18704 0 18760 400
rect 19040 0 19096 400
rect 19376 0 19432 400
rect 19712 0 19768 400
rect 20048 0 20104 400
rect 20384 0 20440 400
rect 20720 0 20776 400
rect 21056 0 21112 400
rect 21392 0 21448 400
rect 21728 0 21784 400
rect 22064 0 22120 400
rect 22400 0 22456 400
rect 22736 0 22792 400
rect 23072 0 23128 400
rect 23408 0 23464 400
rect 23744 0 23800 400
rect 24080 0 24136 400
rect 24416 0 24472 400
rect 24752 0 24808 400
rect 25088 0 25144 400
rect 25424 0 25480 400
rect 25760 0 25816 400
rect 26096 0 26152 400
rect 26432 0 26488 400
rect 26768 0 26824 400
rect 27104 0 27160 400
rect 27440 0 27496 400
rect 27776 0 27832 400
rect 28112 0 28168 400
rect 28448 0 28504 400
rect 28784 0 28840 400
rect 29120 0 29176 400
rect 29456 0 29512 400
rect 29792 0 29848 400
rect 30128 0 30184 400
rect 30464 0 30520 400
rect 30800 0 30856 400
rect 31136 0 31192 400
rect 31472 0 31528 400
rect 31808 0 31864 400
rect 32144 0 32200 400
rect 32480 0 32536 400
rect 32816 0 32872 400
rect 33152 0 33208 400
rect 33488 0 33544 400
rect 33824 0 33880 400
rect 34160 0 34216 400
rect 34496 0 34552 400
rect 34832 0 34888 400
rect 35168 0 35224 400
rect 35504 0 35560 400
rect 35840 0 35896 400
rect 36176 0 36232 400
rect 36512 0 36568 400
rect 36848 0 36904 400
rect 37184 0 37240 400
rect 37520 0 37576 400
rect 37856 0 37912 400
rect 38192 0 38248 400
rect 38528 0 38584 400
rect 38864 0 38920 400
rect 39200 0 39256 400
rect 39536 0 39592 400
rect 39872 0 39928 400
rect 40208 0 40264 400
rect 40544 0 40600 400
rect 40880 0 40936 400
rect 41216 0 41272 400
rect 41552 0 41608 400
rect 41888 0 41944 400
rect 42224 0 42280 400
rect 42560 0 42616 400
rect 42896 0 42952 400
rect 43232 0 43288 400
rect 43568 0 43624 400
rect 43904 0 43960 400
rect 44240 0 44296 400
rect 44576 0 44632 400
rect 44912 0 44968 400
rect 45248 0 45304 400
rect 45584 0 45640 400
rect 45920 0 45976 400
rect 46256 0 46312 400
rect 46592 0 46648 400
rect 46928 0 46984 400
rect 47264 0 47320 400
rect 47600 0 47656 400
rect 47936 0 47992 400
rect 48272 0 48328 400
rect 48608 0 48664 400
rect 48944 0 49000 400
rect 49280 0 49336 400
rect 49616 0 49672 400
rect 49952 0 50008 400
rect 50288 0 50344 400
rect 50624 0 50680 400
rect 50960 0 51016 400
rect 51296 0 51352 400
rect 51632 0 51688 400
rect 51968 0 52024 400
rect 52304 0 52360 400
rect 52640 0 52696 400
rect 52976 0 53032 400
rect 53312 0 53368 400
rect 53648 0 53704 400
rect 53984 0 54040 400
rect 54320 0 54376 400
rect 54656 0 54712 400
rect 54992 0 55048 400
rect 55328 0 55384 400
rect 55664 0 55720 400
rect 56000 0 56056 400
rect 56336 0 56392 400
rect 56672 0 56728 400
rect 57008 0 57064 400
rect 57344 0 57400 400
rect 57680 0 57736 400
rect 58016 0 58072 400
rect 58352 0 58408 400
rect 58688 0 58744 400
rect 59024 0 59080 400
rect 59360 0 59416 400
rect 59696 0 59752 400
rect 60032 0 60088 400
rect 60368 0 60424 400
rect 60704 0 60760 400
rect 61040 0 61096 400
rect 61376 0 61432 400
rect 61712 0 61768 400
rect 62048 0 62104 400
rect 62384 0 62440 400
rect 62720 0 62776 400
rect 63056 0 63112 400
rect 63392 0 63448 400
rect 63728 0 63784 400
rect 64064 0 64120 400
rect 64400 0 64456 400
rect 64736 0 64792 400
rect 65072 0 65128 400
rect 65408 0 65464 400
rect 65744 0 65800 400
rect 66080 0 66136 400
rect 66416 0 66472 400
rect 66752 0 66808 400
rect 67088 0 67144 400
rect 67424 0 67480 400
rect 67760 0 67816 400
rect 68096 0 68152 400
rect 68432 0 68488 400
rect 68768 0 68824 400
rect 69104 0 69160 400
rect 69440 0 69496 400
rect 69776 0 69832 400
rect 70112 0 70168 400
rect 70448 0 70504 400
rect 70784 0 70840 400
rect 71120 0 71176 400
rect 71456 0 71512 400
rect 71792 0 71848 400
rect 72128 0 72184 400
rect 72464 0 72520 400
rect 72800 0 72856 400
rect 73136 0 73192 400
rect 73472 0 73528 400
rect 73808 0 73864 400
rect 74144 0 74200 400
rect 74480 0 74536 400
rect 74816 0 74872 400
rect 75152 0 75208 400
rect 75488 0 75544 400
rect 75824 0 75880 400
rect 76160 0 76216 400
rect 76496 0 76552 400
rect 76832 0 76888 400
rect 77168 0 77224 400
rect 77504 0 77560 400
rect 77840 0 77896 400
rect 78176 0 78232 400
rect 78512 0 78568 400
rect 78848 0 78904 400
rect 79184 0 79240 400
rect 79520 0 79576 400
rect 79856 0 79912 400
rect 80192 0 80248 400
rect 80528 0 80584 400
rect 80864 0 80920 400
rect 81200 0 81256 400
rect 81536 0 81592 400
rect 81872 0 81928 400
rect 82208 0 82264 400
rect 82544 0 82600 400
rect 82880 0 82936 400
rect 83216 0 83272 400
rect 83552 0 83608 400
rect 83888 0 83944 400
rect 84224 0 84280 400
rect 84560 0 84616 400
rect 84896 0 84952 400
rect 85232 0 85288 400
rect 85568 0 85624 400
rect 85904 0 85960 400
rect 86240 0 86296 400
rect 86576 0 86632 400
rect 86912 0 86968 400
rect 87248 0 87304 400
rect 87584 0 87640 400
rect 87920 0 87976 400
rect 88256 0 88312 400
rect 88592 0 88648 400
rect 88928 0 88984 400
rect 89264 0 89320 400
rect 89600 0 89656 400
rect 89936 0 89992 400
rect 90272 0 90328 400
rect 90608 0 90664 400
rect 90944 0 91000 400
rect 91280 0 91336 400
rect 91616 0 91672 400
rect 91952 0 92008 400
rect 92288 0 92344 400
rect 92624 0 92680 400
rect 92960 0 93016 400
rect 93296 0 93352 400
rect 93632 0 93688 400
rect 93968 0 94024 400
rect 94304 0 94360 400
rect 94640 0 94696 400
rect 94976 0 95032 400
rect 95312 0 95368 400
rect 95648 0 95704 400
rect 95984 0 96040 400
rect 96320 0 96376 400
rect 96656 0 96712 400
rect 96992 0 97048 400
rect 97328 0 97384 400
rect 97664 0 97720 400
rect 98000 0 98056 400
rect 98336 0 98392 400
rect 98672 0 98728 400
rect 99008 0 99064 400
rect 99344 0 99400 400
rect 99680 0 99736 400
rect 100016 0 100072 400
rect 100352 0 100408 400
rect 100688 0 100744 400
rect 101024 0 101080 400
rect 101360 0 101416 400
rect 101696 0 101752 400
rect 102032 0 102088 400
rect 102368 0 102424 400
rect 102704 0 102760 400
rect 103040 0 103096 400
rect 103376 0 103432 400
rect 103712 0 103768 400
rect 104048 0 104104 400
rect 104384 0 104440 400
rect 104720 0 104776 400
rect 105056 0 105112 400
rect 105392 0 105448 400
rect 105728 0 105784 400
rect 106064 0 106120 400
rect 106400 0 106456 400
rect 106736 0 106792 400
rect 107072 0 107128 400
rect 107408 0 107464 400
rect 107744 0 107800 400
rect 108080 0 108136 400
rect 108416 0 108472 400
rect 108752 0 108808 400
rect 109088 0 109144 400
rect 109424 0 109480 400
rect 109760 0 109816 400
rect 110096 0 110152 400
rect 110432 0 110488 400
rect 110768 0 110824 400
rect 111104 0 111160 400
rect 111440 0 111496 400
rect 111776 0 111832 400
rect 112112 0 112168 400
rect 112448 0 112504 400
rect 112784 0 112840 400
rect 113120 0 113176 400
rect 113456 0 113512 400
rect 113792 0 113848 400
rect 114128 0 114184 400
rect 114464 0 114520 400
rect 114800 0 114856 400
rect 115136 0 115192 400
rect 115472 0 115528 400
rect 115808 0 115864 400
rect 116144 0 116200 400
rect 116480 0 116536 400
rect 116816 0 116872 400
rect 117152 0 117208 400
rect 117488 0 117544 400
rect 117824 0 117880 400
rect 118160 0 118216 400
rect 118496 0 118552 400
rect 118832 0 118888 400
rect 119168 0 119224 400
rect 119504 0 119560 400
rect 119840 0 119896 400
rect 120176 0 120232 400
rect 120512 0 120568 400
rect 120848 0 120904 400
rect 121184 0 121240 400
rect 121520 0 121576 400
rect 121856 0 121912 400
rect 122192 0 122248 400
rect 122528 0 122584 400
rect 122864 0 122920 400
rect 123200 0 123256 400
rect 123536 0 123592 400
rect 123872 0 123928 400
rect 124208 0 124264 400
rect 124544 0 124600 400
rect 124880 0 124936 400
rect 125216 0 125272 400
rect 125552 0 125608 400
rect 125888 0 125944 400
rect 126224 0 126280 400
rect 126560 0 126616 400
rect 126896 0 126952 400
rect 127232 0 127288 400
rect 127568 0 127624 400
rect 127904 0 127960 400
rect 128240 0 128296 400
rect 128576 0 128632 400
rect 128912 0 128968 400
rect 129248 0 129304 400
rect 129584 0 129640 400
rect 129920 0 129976 400
rect 130256 0 130312 400
rect 130592 0 130648 400
rect 130928 0 130984 400
rect 131264 0 131320 400
rect 131600 0 131656 400
rect 131936 0 131992 400
rect 132272 0 132328 400
rect 132608 0 132664 400
rect 132944 0 133000 400
rect 133280 0 133336 400
rect 133616 0 133672 400
rect 133952 0 134008 400
rect 134288 0 134344 400
rect 134624 0 134680 400
rect 134960 0 135016 400
rect 135296 0 135352 400
rect 135632 0 135688 400
rect 135968 0 136024 400
rect 136304 0 136360 400
rect 136640 0 136696 400
rect 136976 0 137032 400
rect 137312 0 137368 400
rect 137648 0 137704 400
rect 137984 0 138040 400
rect 138320 0 138376 400
rect 138656 0 138712 400
rect 138992 0 139048 400
rect 139328 0 139384 400
rect 139664 0 139720 400
rect 140000 0 140056 400
rect 140336 0 140392 400
rect 140672 0 140728 400
rect 141008 0 141064 400
rect 141344 0 141400 400
rect 141680 0 141736 400
rect 142016 0 142072 400
rect 142352 0 142408 400
rect 142688 0 142744 400
rect 143024 0 143080 400
rect 143360 0 143416 400
rect 143696 0 143752 400
rect 144032 0 144088 400
rect 144368 0 144424 400
rect 144704 0 144760 400
rect 145040 0 145096 400
rect 145376 0 145432 400
rect 145712 0 145768 400
rect 146048 0 146104 400
rect 146384 0 146440 400
rect 146720 0 146776 400
rect 147056 0 147112 400
rect 147392 0 147448 400
rect 147728 0 147784 400
rect 148064 0 148120 400
rect 148400 0 148456 400
rect 148736 0 148792 400
rect 149072 0 149128 400
rect 149408 0 149464 400
rect 149744 0 149800 400
rect 150080 0 150136 400
rect 150416 0 150472 400
rect 150752 0 150808 400
rect 151088 0 151144 400
rect 151424 0 151480 400
rect 151760 0 151816 400
rect 152096 0 152152 400
rect 152432 0 152488 400
rect 152768 0 152824 400
rect 153104 0 153160 400
rect 153440 0 153496 400
rect 153776 0 153832 400
rect 154112 0 154168 400
rect 154448 0 154504 400
rect 154784 0 154840 400
rect 155120 0 155176 400
rect 155456 0 155512 400
rect 155792 0 155848 400
rect 156128 0 156184 400
rect 156464 0 156520 400
rect 156800 0 156856 400
rect 157136 0 157192 400
rect 157472 0 157528 400
rect 157808 0 157864 400
rect 158144 0 158200 400
rect 158480 0 158536 400
rect 158816 0 158872 400
rect 159152 0 159208 400
rect 159488 0 159544 400
rect 159824 0 159880 400
rect 160160 0 160216 400
rect 160496 0 160552 400
rect 160832 0 160888 400
rect 161168 0 161224 400
rect 161504 0 161560 400
rect 161840 0 161896 400
rect 162176 0 162232 400
rect 162512 0 162568 400
rect 162848 0 162904 400
rect 163184 0 163240 400
rect 163520 0 163576 400
rect 163856 0 163912 400
rect 164192 0 164248 400
rect 164528 0 164584 400
rect 164864 0 164920 400
rect 165200 0 165256 400
rect 165536 0 165592 400
rect 165872 0 165928 400
rect 166208 0 166264 400
rect 166544 0 166600 400
rect 166880 0 166936 400
rect 167216 0 167272 400
rect 167552 0 167608 400
rect 167888 0 167944 400
rect 168224 0 168280 400
rect 168560 0 168616 400
rect 168896 0 168952 400
rect 169232 0 169288 400
rect 169568 0 169624 400
rect 169904 0 169960 400
rect 170240 0 170296 400
rect 170576 0 170632 400
rect 170912 0 170968 400
rect 171248 0 171304 400
rect 171584 0 171640 400
rect 171920 0 171976 400
rect 172256 0 172312 400
rect 172592 0 172648 400
rect 172928 0 172984 400
rect 173264 0 173320 400
rect 173600 0 173656 400
rect 173936 0 173992 400
rect 174272 0 174328 400
rect 174608 0 174664 400
rect 174944 0 175000 400
rect 175280 0 175336 400
rect 175616 0 175672 400
rect 175952 0 176008 400
rect 176288 0 176344 400
rect 176624 0 176680 400
rect 176960 0 177016 400
rect 177296 0 177352 400
rect 177632 0 177688 400
rect 177968 0 178024 400
<< obsm2 >>
rect 1638 99570 6746 99783
rect 6862 99570 7362 99783
rect 7478 99570 7978 99783
rect 8094 99570 8594 99783
rect 8710 99570 9210 99783
rect 9326 99570 9826 99783
rect 9942 99570 10442 99783
rect 10558 99570 11058 99783
rect 11174 99570 11674 99783
rect 11790 99570 12290 99783
rect 12406 99570 12906 99783
rect 13022 99570 13522 99783
rect 13638 99570 14138 99783
rect 14254 99570 14754 99783
rect 14870 99570 15370 99783
rect 15486 99570 15986 99783
rect 16102 99570 16602 99783
rect 16718 99570 17218 99783
rect 17334 99570 17834 99783
rect 17950 99570 18450 99783
rect 18566 99570 19066 99783
rect 19182 99570 19682 99783
rect 19798 99570 20298 99783
rect 20414 99570 20914 99783
rect 21030 99570 21530 99783
rect 21646 99570 22146 99783
rect 22262 99570 22762 99783
rect 22878 99570 23378 99783
rect 23494 99570 23994 99783
rect 24110 99570 24610 99783
rect 24726 99570 25226 99783
rect 25342 99570 25842 99783
rect 25958 99570 26458 99783
rect 26574 99570 27074 99783
rect 27190 99570 27690 99783
rect 27806 99570 28306 99783
rect 28422 99570 28922 99783
rect 29038 99570 29538 99783
rect 29654 99570 30154 99783
rect 30270 99570 30770 99783
rect 30886 99570 31386 99783
rect 31502 99570 32002 99783
rect 32118 99570 32618 99783
rect 32734 99570 33234 99783
rect 33350 99570 33850 99783
rect 33966 99570 34466 99783
rect 34582 99570 35082 99783
rect 35198 99570 35698 99783
rect 35814 99570 36314 99783
rect 36430 99570 36930 99783
rect 37046 99570 37546 99783
rect 37662 99570 38162 99783
rect 38278 99570 38778 99783
rect 38894 99570 39394 99783
rect 39510 99570 40010 99783
rect 40126 99570 40626 99783
rect 40742 99570 41242 99783
rect 41358 99570 41858 99783
rect 41974 99570 42474 99783
rect 42590 99570 43090 99783
rect 43206 99570 43706 99783
rect 43822 99570 44322 99783
rect 44438 99570 44938 99783
rect 45054 99570 45554 99783
rect 45670 99570 46170 99783
rect 46286 99570 46786 99783
rect 46902 99570 47402 99783
rect 47518 99570 48018 99783
rect 48134 99570 48634 99783
rect 48750 99570 49250 99783
rect 49366 99570 49866 99783
rect 49982 99570 50482 99783
rect 50598 99570 51098 99783
rect 51214 99570 51714 99783
rect 51830 99570 52330 99783
rect 52446 99570 52946 99783
rect 53062 99570 53562 99783
rect 53678 99570 54178 99783
rect 54294 99570 54794 99783
rect 54910 99570 55410 99783
rect 55526 99570 56026 99783
rect 56142 99570 56642 99783
rect 56758 99570 57258 99783
rect 57374 99570 57874 99783
rect 57990 99570 58490 99783
rect 58606 99570 59106 99783
rect 59222 99570 59722 99783
rect 59838 99570 60338 99783
rect 60454 99570 60954 99783
rect 61070 99570 61570 99783
rect 61686 99570 62186 99783
rect 62302 99570 62802 99783
rect 62918 99570 63418 99783
rect 63534 99570 64034 99783
rect 64150 99570 64650 99783
rect 64766 99570 65266 99783
rect 65382 99570 65882 99783
rect 65998 99570 66498 99783
rect 66614 99570 67114 99783
rect 67230 99570 67730 99783
rect 67846 99570 68346 99783
rect 68462 99570 68962 99783
rect 69078 99570 69578 99783
rect 69694 99570 70194 99783
rect 70310 99570 70810 99783
rect 70926 99570 71426 99783
rect 71542 99570 72042 99783
rect 72158 99570 72658 99783
rect 72774 99570 73274 99783
rect 73390 99570 73890 99783
rect 74006 99570 74506 99783
rect 74622 99570 75122 99783
rect 75238 99570 75738 99783
rect 75854 99570 76354 99783
rect 76470 99570 76970 99783
rect 77086 99570 77586 99783
rect 77702 99570 78202 99783
rect 78318 99570 78818 99783
rect 78934 99570 79434 99783
rect 79550 99570 80050 99783
rect 80166 99570 80666 99783
rect 80782 99570 81282 99783
rect 81398 99570 81898 99783
rect 82014 99570 82514 99783
rect 82630 99570 83130 99783
rect 83246 99570 83746 99783
rect 83862 99570 84362 99783
rect 84478 99570 84978 99783
rect 85094 99570 85594 99783
rect 85710 99570 86210 99783
rect 86326 99570 86826 99783
rect 86942 99570 87442 99783
rect 87558 99570 88058 99783
rect 88174 99570 88674 99783
rect 88790 99570 89290 99783
rect 89406 99570 89906 99783
rect 90022 99570 90522 99783
rect 90638 99570 91138 99783
rect 91254 99570 91754 99783
rect 91870 99570 92370 99783
rect 92486 99570 92986 99783
rect 93102 99570 93602 99783
rect 93718 99570 94218 99783
rect 94334 99570 94834 99783
rect 94950 99570 95450 99783
rect 95566 99570 96066 99783
rect 96182 99570 96682 99783
rect 96798 99570 97298 99783
rect 97414 99570 97914 99783
rect 98030 99570 98530 99783
rect 98646 99570 99146 99783
rect 99262 99570 99762 99783
rect 99878 99570 100378 99783
rect 100494 99570 100994 99783
rect 101110 99570 101610 99783
rect 101726 99570 102226 99783
rect 102342 99570 102842 99783
rect 102958 99570 103458 99783
rect 103574 99570 104074 99783
rect 104190 99570 104690 99783
rect 104806 99570 105306 99783
rect 105422 99570 105922 99783
rect 106038 99570 106538 99783
rect 106654 99570 107154 99783
rect 107270 99570 107770 99783
rect 107886 99570 108386 99783
rect 108502 99570 109002 99783
rect 109118 99570 109618 99783
rect 109734 99570 110234 99783
rect 110350 99570 110850 99783
rect 110966 99570 111466 99783
rect 111582 99570 112082 99783
rect 112198 99570 112698 99783
rect 112814 99570 113314 99783
rect 113430 99570 113930 99783
rect 114046 99570 114546 99783
rect 114662 99570 115162 99783
rect 115278 99570 115778 99783
rect 115894 99570 116394 99783
rect 116510 99570 117010 99783
rect 117126 99570 117626 99783
rect 117742 99570 118242 99783
rect 118358 99570 118858 99783
rect 118974 99570 119474 99783
rect 119590 99570 120090 99783
rect 120206 99570 120706 99783
rect 120822 99570 121322 99783
rect 121438 99570 121938 99783
rect 122054 99570 122554 99783
rect 122670 99570 123170 99783
rect 123286 99570 123786 99783
rect 123902 99570 124402 99783
rect 124518 99570 125018 99783
rect 125134 99570 125634 99783
rect 125750 99570 126250 99783
rect 126366 99570 126866 99783
rect 126982 99570 127482 99783
rect 127598 99570 128098 99783
rect 128214 99570 128714 99783
rect 128830 99570 129330 99783
rect 129446 99570 129946 99783
rect 130062 99570 130562 99783
rect 130678 99570 131178 99783
rect 131294 99570 131794 99783
rect 131910 99570 132410 99783
rect 132526 99570 133026 99783
rect 133142 99570 133642 99783
rect 133758 99570 134258 99783
rect 134374 99570 134874 99783
rect 134990 99570 135490 99783
rect 135606 99570 136106 99783
rect 136222 99570 136722 99783
rect 136838 99570 137338 99783
rect 137454 99570 137954 99783
rect 138070 99570 138570 99783
rect 138686 99570 139186 99783
rect 139302 99570 139802 99783
rect 139918 99570 140418 99783
rect 140534 99570 141034 99783
rect 141150 99570 141650 99783
rect 141766 99570 142266 99783
rect 142382 99570 142882 99783
rect 142998 99570 143498 99783
rect 143614 99570 144114 99783
rect 144230 99570 144730 99783
rect 144846 99570 145346 99783
rect 145462 99570 145962 99783
rect 146078 99570 146578 99783
rect 146694 99570 147194 99783
rect 147310 99570 147810 99783
rect 147926 99570 148426 99783
rect 148542 99570 149042 99783
rect 149158 99570 149658 99783
rect 149774 99570 150274 99783
rect 150390 99570 150890 99783
rect 151006 99570 151506 99783
rect 151622 99570 152122 99783
rect 152238 99570 152738 99783
rect 152854 99570 153354 99783
rect 153470 99570 153970 99783
rect 154086 99570 154586 99783
rect 154702 99570 155202 99783
rect 155318 99570 155818 99783
rect 155934 99570 156434 99783
rect 156550 99570 157050 99783
rect 157166 99570 157666 99783
rect 157782 99570 158282 99783
rect 158398 99570 158898 99783
rect 159014 99570 159514 99783
rect 159630 99570 160130 99783
rect 160246 99570 160746 99783
rect 160862 99570 161362 99783
rect 161478 99570 161978 99783
rect 162094 99570 162594 99783
rect 162710 99570 163210 99783
rect 163326 99570 163826 99783
rect 163942 99570 164442 99783
rect 164558 99570 165058 99783
rect 165174 99570 165674 99783
rect 165790 99570 166290 99783
rect 166406 99570 166906 99783
rect 167022 99570 167522 99783
rect 167638 99570 168138 99783
rect 168254 99570 168754 99783
rect 168870 99570 169370 99783
rect 169486 99570 169986 99783
rect 170102 99570 170602 99783
rect 170718 99570 171218 99783
rect 171334 99570 171834 99783
rect 171950 99570 172450 99783
rect 172566 99570 173066 99783
rect 173182 99570 179074 99783
rect 1638 430 179074 99570
rect 1638 9 1874 430
rect 1990 9 2210 430
rect 2326 9 2546 430
rect 2662 9 2882 430
rect 2998 9 3218 430
rect 3334 9 3554 430
rect 3670 9 3890 430
rect 4006 9 4226 430
rect 4342 9 4562 430
rect 4678 9 4898 430
rect 5014 9 5234 430
rect 5350 9 5570 430
rect 5686 9 5906 430
rect 6022 9 6242 430
rect 6358 9 6578 430
rect 6694 9 6914 430
rect 7030 9 7250 430
rect 7366 9 7586 430
rect 7702 9 7922 430
rect 8038 9 8258 430
rect 8374 9 8594 430
rect 8710 9 8930 430
rect 9046 9 9266 430
rect 9382 9 9602 430
rect 9718 9 9938 430
rect 10054 9 10274 430
rect 10390 9 10610 430
rect 10726 9 10946 430
rect 11062 9 11282 430
rect 11398 9 11618 430
rect 11734 9 11954 430
rect 12070 9 12290 430
rect 12406 9 12626 430
rect 12742 9 12962 430
rect 13078 9 13298 430
rect 13414 9 13634 430
rect 13750 9 13970 430
rect 14086 9 14306 430
rect 14422 9 14642 430
rect 14758 9 14978 430
rect 15094 9 15314 430
rect 15430 9 15650 430
rect 15766 9 15986 430
rect 16102 9 16322 430
rect 16438 9 16658 430
rect 16774 9 16994 430
rect 17110 9 17330 430
rect 17446 9 17666 430
rect 17782 9 18002 430
rect 18118 9 18338 430
rect 18454 9 18674 430
rect 18790 9 19010 430
rect 19126 9 19346 430
rect 19462 9 19682 430
rect 19798 9 20018 430
rect 20134 9 20354 430
rect 20470 9 20690 430
rect 20806 9 21026 430
rect 21142 9 21362 430
rect 21478 9 21698 430
rect 21814 9 22034 430
rect 22150 9 22370 430
rect 22486 9 22706 430
rect 22822 9 23042 430
rect 23158 9 23378 430
rect 23494 9 23714 430
rect 23830 9 24050 430
rect 24166 9 24386 430
rect 24502 9 24722 430
rect 24838 9 25058 430
rect 25174 9 25394 430
rect 25510 9 25730 430
rect 25846 9 26066 430
rect 26182 9 26402 430
rect 26518 9 26738 430
rect 26854 9 27074 430
rect 27190 9 27410 430
rect 27526 9 27746 430
rect 27862 9 28082 430
rect 28198 9 28418 430
rect 28534 9 28754 430
rect 28870 9 29090 430
rect 29206 9 29426 430
rect 29542 9 29762 430
rect 29878 9 30098 430
rect 30214 9 30434 430
rect 30550 9 30770 430
rect 30886 9 31106 430
rect 31222 9 31442 430
rect 31558 9 31778 430
rect 31894 9 32114 430
rect 32230 9 32450 430
rect 32566 9 32786 430
rect 32902 9 33122 430
rect 33238 9 33458 430
rect 33574 9 33794 430
rect 33910 9 34130 430
rect 34246 9 34466 430
rect 34582 9 34802 430
rect 34918 9 35138 430
rect 35254 9 35474 430
rect 35590 9 35810 430
rect 35926 9 36146 430
rect 36262 9 36482 430
rect 36598 9 36818 430
rect 36934 9 37154 430
rect 37270 9 37490 430
rect 37606 9 37826 430
rect 37942 9 38162 430
rect 38278 9 38498 430
rect 38614 9 38834 430
rect 38950 9 39170 430
rect 39286 9 39506 430
rect 39622 9 39842 430
rect 39958 9 40178 430
rect 40294 9 40514 430
rect 40630 9 40850 430
rect 40966 9 41186 430
rect 41302 9 41522 430
rect 41638 9 41858 430
rect 41974 9 42194 430
rect 42310 9 42530 430
rect 42646 9 42866 430
rect 42982 9 43202 430
rect 43318 9 43538 430
rect 43654 9 43874 430
rect 43990 9 44210 430
rect 44326 9 44546 430
rect 44662 9 44882 430
rect 44998 9 45218 430
rect 45334 9 45554 430
rect 45670 9 45890 430
rect 46006 9 46226 430
rect 46342 9 46562 430
rect 46678 9 46898 430
rect 47014 9 47234 430
rect 47350 9 47570 430
rect 47686 9 47906 430
rect 48022 9 48242 430
rect 48358 9 48578 430
rect 48694 9 48914 430
rect 49030 9 49250 430
rect 49366 9 49586 430
rect 49702 9 49922 430
rect 50038 9 50258 430
rect 50374 9 50594 430
rect 50710 9 50930 430
rect 51046 9 51266 430
rect 51382 9 51602 430
rect 51718 9 51938 430
rect 52054 9 52274 430
rect 52390 9 52610 430
rect 52726 9 52946 430
rect 53062 9 53282 430
rect 53398 9 53618 430
rect 53734 9 53954 430
rect 54070 9 54290 430
rect 54406 9 54626 430
rect 54742 9 54962 430
rect 55078 9 55298 430
rect 55414 9 55634 430
rect 55750 9 55970 430
rect 56086 9 56306 430
rect 56422 9 56642 430
rect 56758 9 56978 430
rect 57094 9 57314 430
rect 57430 9 57650 430
rect 57766 9 57986 430
rect 58102 9 58322 430
rect 58438 9 58658 430
rect 58774 9 58994 430
rect 59110 9 59330 430
rect 59446 9 59666 430
rect 59782 9 60002 430
rect 60118 9 60338 430
rect 60454 9 60674 430
rect 60790 9 61010 430
rect 61126 9 61346 430
rect 61462 9 61682 430
rect 61798 9 62018 430
rect 62134 9 62354 430
rect 62470 9 62690 430
rect 62806 9 63026 430
rect 63142 9 63362 430
rect 63478 9 63698 430
rect 63814 9 64034 430
rect 64150 9 64370 430
rect 64486 9 64706 430
rect 64822 9 65042 430
rect 65158 9 65378 430
rect 65494 9 65714 430
rect 65830 9 66050 430
rect 66166 9 66386 430
rect 66502 9 66722 430
rect 66838 9 67058 430
rect 67174 9 67394 430
rect 67510 9 67730 430
rect 67846 9 68066 430
rect 68182 9 68402 430
rect 68518 9 68738 430
rect 68854 9 69074 430
rect 69190 9 69410 430
rect 69526 9 69746 430
rect 69862 9 70082 430
rect 70198 9 70418 430
rect 70534 9 70754 430
rect 70870 9 71090 430
rect 71206 9 71426 430
rect 71542 9 71762 430
rect 71878 9 72098 430
rect 72214 9 72434 430
rect 72550 9 72770 430
rect 72886 9 73106 430
rect 73222 9 73442 430
rect 73558 9 73778 430
rect 73894 9 74114 430
rect 74230 9 74450 430
rect 74566 9 74786 430
rect 74902 9 75122 430
rect 75238 9 75458 430
rect 75574 9 75794 430
rect 75910 9 76130 430
rect 76246 9 76466 430
rect 76582 9 76802 430
rect 76918 9 77138 430
rect 77254 9 77474 430
rect 77590 9 77810 430
rect 77926 9 78146 430
rect 78262 9 78482 430
rect 78598 9 78818 430
rect 78934 9 79154 430
rect 79270 9 79490 430
rect 79606 9 79826 430
rect 79942 9 80162 430
rect 80278 9 80498 430
rect 80614 9 80834 430
rect 80950 9 81170 430
rect 81286 9 81506 430
rect 81622 9 81842 430
rect 81958 9 82178 430
rect 82294 9 82514 430
rect 82630 9 82850 430
rect 82966 9 83186 430
rect 83302 9 83522 430
rect 83638 9 83858 430
rect 83974 9 84194 430
rect 84310 9 84530 430
rect 84646 9 84866 430
rect 84982 9 85202 430
rect 85318 9 85538 430
rect 85654 9 85874 430
rect 85990 9 86210 430
rect 86326 9 86546 430
rect 86662 9 86882 430
rect 86998 9 87218 430
rect 87334 9 87554 430
rect 87670 9 87890 430
rect 88006 9 88226 430
rect 88342 9 88562 430
rect 88678 9 88898 430
rect 89014 9 89234 430
rect 89350 9 89570 430
rect 89686 9 89906 430
rect 90022 9 90242 430
rect 90358 9 90578 430
rect 90694 9 90914 430
rect 91030 9 91250 430
rect 91366 9 91586 430
rect 91702 9 91922 430
rect 92038 9 92258 430
rect 92374 9 92594 430
rect 92710 9 92930 430
rect 93046 9 93266 430
rect 93382 9 93602 430
rect 93718 9 93938 430
rect 94054 9 94274 430
rect 94390 9 94610 430
rect 94726 9 94946 430
rect 95062 9 95282 430
rect 95398 9 95618 430
rect 95734 9 95954 430
rect 96070 9 96290 430
rect 96406 9 96626 430
rect 96742 9 96962 430
rect 97078 9 97298 430
rect 97414 9 97634 430
rect 97750 9 97970 430
rect 98086 9 98306 430
rect 98422 9 98642 430
rect 98758 9 98978 430
rect 99094 9 99314 430
rect 99430 9 99650 430
rect 99766 9 99986 430
rect 100102 9 100322 430
rect 100438 9 100658 430
rect 100774 9 100994 430
rect 101110 9 101330 430
rect 101446 9 101666 430
rect 101782 9 102002 430
rect 102118 9 102338 430
rect 102454 9 102674 430
rect 102790 9 103010 430
rect 103126 9 103346 430
rect 103462 9 103682 430
rect 103798 9 104018 430
rect 104134 9 104354 430
rect 104470 9 104690 430
rect 104806 9 105026 430
rect 105142 9 105362 430
rect 105478 9 105698 430
rect 105814 9 106034 430
rect 106150 9 106370 430
rect 106486 9 106706 430
rect 106822 9 107042 430
rect 107158 9 107378 430
rect 107494 9 107714 430
rect 107830 9 108050 430
rect 108166 9 108386 430
rect 108502 9 108722 430
rect 108838 9 109058 430
rect 109174 9 109394 430
rect 109510 9 109730 430
rect 109846 9 110066 430
rect 110182 9 110402 430
rect 110518 9 110738 430
rect 110854 9 111074 430
rect 111190 9 111410 430
rect 111526 9 111746 430
rect 111862 9 112082 430
rect 112198 9 112418 430
rect 112534 9 112754 430
rect 112870 9 113090 430
rect 113206 9 113426 430
rect 113542 9 113762 430
rect 113878 9 114098 430
rect 114214 9 114434 430
rect 114550 9 114770 430
rect 114886 9 115106 430
rect 115222 9 115442 430
rect 115558 9 115778 430
rect 115894 9 116114 430
rect 116230 9 116450 430
rect 116566 9 116786 430
rect 116902 9 117122 430
rect 117238 9 117458 430
rect 117574 9 117794 430
rect 117910 9 118130 430
rect 118246 9 118466 430
rect 118582 9 118802 430
rect 118918 9 119138 430
rect 119254 9 119474 430
rect 119590 9 119810 430
rect 119926 9 120146 430
rect 120262 9 120482 430
rect 120598 9 120818 430
rect 120934 9 121154 430
rect 121270 9 121490 430
rect 121606 9 121826 430
rect 121942 9 122162 430
rect 122278 9 122498 430
rect 122614 9 122834 430
rect 122950 9 123170 430
rect 123286 9 123506 430
rect 123622 9 123842 430
rect 123958 9 124178 430
rect 124294 9 124514 430
rect 124630 9 124850 430
rect 124966 9 125186 430
rect 125302 9 125522 430
rect 125638 9 125858 430
rect 125974 9 126194 430
rect 126310 9 126530 430
rect 126646 9 126866 430
rect 126982 9 127202 430
rect 127318 9 127538 430
rect 127654 9 127874 430
rect 127990 9 128210 430
rect 128326 9 128546 430
rect 128662 9 128882 430
rect 128998 9 129218 430
rect 129334 9 129554 430
rect 129670 9 129890 430
rect 130006 9 130226 430
rect 130342 9 130562 430
rect 130678 9 130898 430
rect 131014 9 131234 430
rect 131350 9 131570 430
rect 131686 9 131906 430
rect 132022 9 132242 430
rect 132358 9 132578 430
rect 132694 9 132914 430
rect 133030 9 133250 430
rect 133366 9 133586 430
rect 133702 9 133922 430
rect 134038 9 134258 430
rect 134374 9 134594 430
rect 134710 9 134930 430
rect 135046 9 135266 430
rect 135382 9 135602 430
rect 135718 9 135938 430
rect 136054 9 136274 430
rect 136390 9 136610 430
rect 136726 9 136946 430
rect 137062 9 137282 430
rect 137398 9 137618 430
rect 137734 9 137954 430
rect 138070 9 138290 430
rect 138406 9 138626 430
rect 138742 9 138962 430
rect 139078 9 139298 430
rect 139414 9 139634 430
rect 139750 9 139970 430
rect 140086 9 140306 430
rect 140422 9 140642 430
rect 140758 9 140978 430
rect 141094 9 141314 430
rect 141430 9 141650 430
rect 141766 9 141986 430
rect 142102 9 142322 430
rect 142438 9 142658 430
rect 142774 9 142994 430
rect 143110 9 143330 430
rect 143446 9 143666 430
rect 143782 9 144002 430
rect 144118 9 144338 430
rect 144454 9 144674 430
rect 144790 9 145010 430
rect 145126 9 145346 430
rect 145462 9 145682 430
rect 145798 9 146018 430
rect 146134 9 146354 430
rect 146470 9 146690 430
rect 146806 9 147026 430
rect 147142 9 147362 430
rect 147478 9 147698 430
rect 147814 9 148034 430
rect 148150 9 148370 430
rect 148486 9 148706 430
rect 148822 9 149042 430
rect 149158 9 149378 430
rect 149494 9 149714 430
rect 149830 9 150050 430
rect 150166 9 150386 430
rect 150502 9 150722 430
rect 150838 9 151058 430
rect 151174 9 151394 430
rect 151510 9 151730 430
rect 151846 9 152066 430
rect 152182 9 152402 430
rect 152518 9 152738 430
rect 152854 9 153074 430
rect 153190 9 153410 430
rect 153526 9 153746 430
rect 153862 9 154082 430
rect 154198 9 154418 430
rect 154534 9 154754 430
rect 154870 9 155090 430
rect 155206 9 155426 430
rect 155542 9 155762 430
rect 155878 9 156098 430
rect 156214 9 156434 430
rect 156550 9 156770 430
rect 156886 9 157106 430
rect 157222 9 157442 430
rect 157558 9 157778 430
rect 157894 9 158114 430
rect 158230 9 158450 430
rect 158566 9 158786 430
rect 158902 9 159122 430
rect 159238 9 159458 430
rect 159574 9 159794 430
rect 159910 9 160130 430
rect 160246 9 160466 430
rect 160582 9 160802 430
rect 160918 9 161138 430
rect 161254 9 161474 430
rect 161590 9 161810 430
rect 161926 9 162146 430
rect 162262 9 162482 430
rect 162598 9 162818 430
rect 162934 9 163154 430
rect 163270 9 163490 430
rect 163606 9 163826 430
rect 163942 9 164162 430
rect 164278 9 164498 430
rect 164614 9 164834 430
rect 164950 9 165170 430
rect 165286 9 165506 430
rect 165622 9 165842 430
rect 165958 9 166178 430
rect 166294 9 166514 430
rect 166630 9 166850 430
rect 166966 9 167186 430
rect 167302 9 167522 430
rect 167638 9 167858 430
rect 167974 9 168194 430
rect 168310 9 168530 430
rect 168646 9 168866 430
rect 168982 9 169202 430
rect 169318 9 169538 430
rect 169654 9 169874 430
rect 169990 9 170210 430
rect 170326 9 170546 430
rect 170662 9 170882 430
rect 170998 9 171218 430
rect 171334 9 171554 430
rect 171670 9 171890 430
rect 172006 9 172226 430
rect 172342 9 172562 430
rect 172678 9 172898 430
rect 173014 9 173234 430
rect 173350 9 173570 430
rect 173686 9 173906 430
rect 174022 9 174242 430
rect 174358 9 174578 430
rect 174694 9 174914 430
rect 175030 9 175250 430
rect 175366 9 175586 430
rect 175702 9 175922 430
rect 176038 9 176258 430
rect 176374 9 176594 430
rect 176710 9 176930 430
rect 177046 9 177266 430
rect 177382 9 177602 430
rect 177718 9 177938 430
rect 178054 9 179074 430
<< obsm3 >>
rect 1633 14 179079 99778
<< metal4 >>
rect 2224 1538 2384 98422
rect 9904 1538 10064 98422
rect 17584 1538 17744 98422
rect 25264 1538 25424 98422
rect 32944 1538 33104 98422
rect 40624 1538 40784 98422
rect 48304 1538 48464 98422
rect 55984 1538 56144 98422
rect 63664 1538 63824 98422
rect 71344 1538 71504 98422
rect 79024 1538 79184 98422
rect 86704 1538 86864 98422
rect 94384 1538 94544 98422
rect 102064 1538 102224 98422
rect 109744 1538 109904 98422
rect 117424 1538 117584 98422
rect 125104 1538 125264 98422
rect 132784 1538 132944 98422
rect 140464 1538 140624 98422
rect 148144 1538 148304 98422
rect 155824 1538 155984 98422
rect 163504 1538 163664 98422
rect 171184 1538 171344 98422
rect 178864 1538 179024 98422
<< obsm4 >>
rect 15974 98452 137690 99447
rect 15974 2641 17554 98452
rect 17774 2641 25234 98452
rect 25454 2641 32914 98452
rect 33134 2641 40594 98452
rect 40814 2641 48274 98452
rect 48494 2641 55954 98452
rect 56174 2641 63634 98452
rect 63854 2641 71314 98452
rect 71534 2641 78994 98452
rect 79214 2641 86674 98452
rect 86894 2641 94354 98452
rect 94574 2641 102034 98452
rect 102254 2641 109714 98452
rect 109934 2641 117394 98452
rect 117614 2641 125074 98452
rect 125294 2641 132754 98452
rect 132974 2641 137690 98452
<< labels >>
rlabel metal2 s 172480 99600 172536 100000 6 Serial_input
port 1 nsew signal input
rlabel metal2 s 173096 99600 173152 100000 6 Serial_output
port 2 nsew signal output
rlabel metal2 s 166544 0 166600 400 6 analog_io[0]
port 3 nsew signal bidirectional
rlabel metal2 s 169904 0 169960 400 6 analog_io[10]
port 4 nsew signal bidirectional
rlabel metal2 s 170240 0 170296 400 6 analog_io[11]
port 5 nsew signal bidirectional
rlabel metal2 s 170576 0 170632 400 6 analog_io[12]
port 6 nsew signal bidirectional
rlabel metal2 s 170912 0 170968 400 6 analog_io[13]
port 7 nsew signal bidirectional
rlabel metal2 s 171248 0 171304 400 6 analog_io[14]
port 8 nsew signal bidirectional
rlabel metal2 s 171584 0 171640 400 6 analog_io[15]
port 9 nsew signal bidirectional
rlabel metal2 s 171920 0 171976 400 6 analog_io[16]
port 10 nsew signal bidirectional
rlabel metal2 s 172256 0 172312 400 6 analog_io[17]
port 11 nsew signal bidirectional
rlabel metal2 s 172592 0 172648 400 6 analog_io[18]
port 12 nsew signal bidirectional
rlabel metal2 s 172928 0 172984 400 6 analog_io[19]
port 13 nsew signal bidirectional
rlabel metal2 s 166880 0 166936 400 6 analog_io[1]
port 14 nsew signal bidirectional
rlabel metal2 s 173264 0 173320 400 6 analog_io[20]
port 15 nsew signal bidirectional
rlabel metal2 s 173600 0 173656 400 6 analog_io[21]
port 16 nsew signal bidirectional
rlabel metal2 s 173936 0 173992 400 6 analog_io[22]
port 17 nsew signal bidirectional
rlabel metal2 s 174272 0 174328 400 6 analog_io[23]
port 18 nsew signal bidirectional
rlabel metal2 s 174608 0 174664 400 6 analog_io[24]
port 19 nsew signal bidirectional
rlabel metal2 s 174944 0 175000 400 6 analog_io[25]
port 20 nsew signal bidirectional
rlabel metal2 s 175280 0 175336 400 6 analog_io[26]
port 21 nsew signal bidirectional
rlabel metal2 s 175616 0 175672 400 6 analog_io[27]
port 22 nsew signal bidirectional
rlabel metal2 s 175952 0 176008 400 6 analog_io[28]
port 23 nsew signal bidirectional
rlabel metal2 s 167216 0 167272 400 6 analog_io[2]
port 24 nsew signal bidirectional
rlabel metal2 s 167552 0 167608 400 6 analog_io[3]
port 25 nsew signal bidirectional
rlabel metal2 s 167888 0 167944 400 6 analog_io[4]
port 26 nsew signal bidirectional
rlabel metal2 s 168224 0 168280 400 6 analog_io[5]
port 27 nsew signal bidirectional
rlabel metal2 s 168560 0 168616 400 6 analog_io[6]
port 28 nsew signal bidirectional
rlabel metal2 s 168896 0 168952 400 6 analog_io[7]
port 29 nsew signal bidirectional
rlabel metal2 s 169232 0 169288 400 6 analog_io[8]
port 30 nsew signal bidirectional
rlabel metal2 s 169568 0 169624 400 6 analog_io[9]
port 31 nsew signal bidirectional
rlabel metal2 s 177296 0 177352 400 6 clk
port 32 nsew signal output
rlabel metal2 s 111496 99600 111552 100000 6 data_mem_addr[0]
port 33 nsew signal output
rlabel metal2 s 113960 99600 114016 100000 6 data_mem_addr[1]
port 34 nsew signal output
rlabel metal2 s 116424 99600 116480 100000 6 data_mem_addr[2]
port 35 nsew signal output
rlabel metal2 s 118888 99600 118944 100000 6 data_mem_addr[3]
port 36 nsew signal output
rlabel metal2 s 121352 99600 121408 100000 6 data_mem_addr[4]
port 37 nsew signal output
rlabel metal2 s 123816 99600 123872 100000 6 data_mem_addr[5]
port 38 nsew signal output
rlabel metal2 s 126280 99600 126336 100000 6 data_mem_addr[6]
port 39 nsew signal output
rlabel metal2 s 128744 99600 128800 100000 6 data_mem_addr[7]
port 40 nsew signal output
rlabel metal2 s 110264 99600 110320 100000 6 data_mem_sel
port 41 nsew signal output
rlabel metal2 s 112112 99600 112168 100000 6 data_read_data[0]
port 42 nsew signal input
rlabel metal2 s 133672 99600 133728 100000 6 data_read_data[10]
port 43 nsew signal input
rlabel metal2 s 134904 99600 134960 100000 6 data_read_data[11]
port 44 nsew signal input
rlabel metal2 s 136136 99600 136192 100000 6 data_read_data[12]
port 45 nsew signal input
rlabel metal2 s 137368 99600 137424 100000 6 data_read_data[13]
port 46 nsew signal input
rlabel metal2 s 138600 99600 138656 100000 6 data_read_data[14]
port 47 nsew signal input
rlabel metal2 s 139832 99600 139888 100000 6 data_read_data[15]
port 48 nsew signal input
rlabel metal2 s 114576 99600 114632 100000 6 data_read_data[1]
port 49 nsew signal input
rlabel metal2 s 117040 99600 117096 100000 6 data_read_data[2]
port 50 nsew signal input
rlabel metal2 s 119504 99600 119560 100000 6 data_read_data[3]
port 51 nsew signal input
rlabel metal2 s 121968 99600 122024 100000 6 data_read_data[4]
port 52 nsew signal input
rlabel metal2 s 124432 99600 124488 100000 6 data_read_data[5]
port 53 nsew signal input
rlabel metal2 s 126896 99600 126952 100000 6 data_read_data[6]
port 54 nsew signal input
rlabel metal2 s 129360 99600 129416 100000 6 data_read_data[7]
port 55 nsew signal input
rlabel metal2 s 131208 99600 131264 100000 6 data_read_data[8]
port 56 nsew signal input
rlabel metal2 s 132440 99600 132496 100000 6 data_read_data[9]
port 57 nsew signal input
rlabel metal2 s 112728 99600 112784 100000 6 data_write_data[0]
port 58 nsew signal output
rlabel metal2 s 134288 99600 134344 100000 6 data_write_data[10]
port 59 nsew signal output
rlabel metal2 s 135520 99600 135576 100000 6 data_write_data[11]
port 60 nsew signal output
rlabel metal2 s 136752 99600 136808 100000 6 data_write_data[12]
port 61 nsew signal output
rlabel metal2 s 137984 99600 138040 100000 6 data_write_data[13]
port 62 nsew signal output
rlabel metal2 s 139216 99600 139272 100000 6 data_write_data[14]
port 63 nsew signal output
rlabel metal2 s 140448 99600 140504 100000 6 data_write_data[15]
port 64 nsew signal output
rlabel metal2 s 115192 99600 115248 100000 6 data_write_data[1]
port 65 nsew signal output
rlabel metal2 s 117656 99600 117712 100000 6 data_write_data[2]
port 66 nsew signal output
rlabel metal2 s 120120 99600 120176 100000 6 data_write_data[3]
port 67 nsew signal output
rlabel metal2 s 122584 99600 122640 100000 6 data_write_data[4]
port 68 nsew signal output
rlabel metal2 s 125048 99600 125104 100000 6 data_write_data[5]
port 69 nsew signal output
rlabel metal2 s 127512 99600 127568 100000 6 data_write_data[6]
port 70 nsew signal output
rlabel metal2 s 129976 99600 130032 100000 6 data_write_data[7]
port 71 nsew signal output
rlabel metal2 s 131824 99600 131880 100000 6 data_write_data[8]
port 72 nsew signal output
rlabel metal2 s 133056 99600 133112 100000 6 data_write_data[9]
port 73 nsew signal output
rlabel metal2 s 110880 99600 110936 100000 6 dataw_en
port 74 nsew signal output
rlabel metal2 s 113344 99600 113400 100000 6 dataw_en_8bit[0]
port 75 nsew signal output
rlabel metal2 s 115808 99600 115864 100000 6 dataw_en_8bit[1]
port 76 nsew signal output
rlabel metal2 s 118272 99600 118328 100000 6 dataw_en_8bit[2]
port 77 nsew signal output
rlabel metal2 s 120736 99600 120792 100000 6 dataw_en_8bit[3]
port 78 nsew signal output
rlabel metal2 s 123200 99600 123256 100000 6 dataw_en_8bit[4]
port 79 nsew signal output
rlabel metal2 s 125664 99600 125720 100000 6 dataw_en_8bit[5]
port 80 nsew signal output
rlabel metal2 s 128128 99600 128184 100000 6 dataw_en_8bit[6]
port 81 nsew signal output
rlabel metal2 s 130592 99600 130648 100000 6 dataw_en_8bit[7]
port 82 nsew signal output
rlabel metal2 s 171864 99600 171920 100000 6 hlt
port 83 nsew signal input
rlabel metal2 s 142296 99600 142352 100000 6 instr[0]
port 84 nsew signal input
rlabel metal2 s 164472 99600 164528 100000 6 instr[10]
port 85 nsew signal input
rlabel metal2 s 165704 99600 165760 100000 6 instr[11]
port 86 nsew signal input
rlabel metal2 s 166936 99600 166992 100000 6 instr[12]
port 87 nsew signal input
rlabel metal2 s 168168 99600 168224 100000 6 instr[13]
port 88 nsew signal input
rlabel metal2 s 169400 99600 169456 100000 6 instr[14]
port 89 nsew signal input
rlabel metal2 s 170632 99600 170688 100000 6 instr[15]
port 90 nsew signal input
rlabel metal2 s 144760 99600 144816 100000 6 instr[1]
port 91 nsew signal input
rlabel metal2 s 147224 99600 147280 100000 6 instr[2]
port 92 nsew signal input
rlabel metal2 s 149688 99600 149744 100000 6 instr[3]
port 93 nsew signal input
rlabel metal2 s 152152 99600 152208 100000 6 instr[4]
port 94 nsew signal input
rlabel metal2 s 154616 99600 154672 100000 6 instr[5]
port 95 nsew signal input
rlabel metal2 s 157080 99600 157136 100000 6 instr[6]
port 96 nsew signal input
rlabel metal2 s 159544 99600 159600 100000 6 instr[7]
port 97 nsew signal input
rlabel metal2 s 162008 99600 162064 100000 6 instr[8]
port 98 nsew signal input
rlabel metal2 s 163240 99600 163296 100000 6 instr[9]
port 99 nsew signal input
rlabel metal2 s 142912 99600 142968 100000 6 instr_mem_addr[0]
port 100 nsew signal output
rlabel metal2 s 145376 99600 145432 100000 6 instr_mem_addr[1]
port 101 nsew signal output
rlabel metal2 s 147840 99600 147896 100000 6 instr_mem_addr[2]
port 102 nsew signal output
rlabel metal2 s 150304 99600 150360 100000 6 instr_mem_addr[3]
port 103 nsew signal output
rlabel metal2 s 152768 99600 152824 100000 6 instr_mem_addr[4]
port 104 nsew signal output
rlabel metal2 s 155232 99600 155288 100000 6 instr_mem_addr[5]
port 105 nsew signal output
rlabel metal2 s 157696 99600 157752 100000 6 instr_mem_addr[6]
port 106 nsew signal output
rlabel metal2 s 160160 99600 160216 100000 6 instr_mem_addr[7]
port 107 nsew signal output
rlabel metal2 s 141064 99600 141120 100000 6 instr_mem_sel
port 108 nsew signal output
rlabel metal2 s 143528 99600 143584 100000 6 instr_write_data[0]
port 109 nsew signal output
rlabel metal2 s 165088 99600 165144 100000 6 instr_write_data[10]
port 110 nsew signal output
rlabel metal2 s 166320 99600 166376 100000 6 instr_write_data[11]
port 111 nsew signal output
rlabel metal2 s 167552 99600 167608 100000 6 instr_write_data[12]
port 112 nsew signal output
rlabel metal2 s 168784 99600 168840 100000 6 instr_write_data[13]
port 113 nsew signal output
rlabel metal2 s 170016 99600 170072 100000 6 instr_write_data[14]
port 114 nsew signal output
rlabel metal2 s 171248 99600 171304 100000 6 instr_write_data[15]
port 115 nsew signal output
rlabel metal2 s 145992 99600 146048 100000 6 instr_write_data[1]
port 116 nsew signal output
rlabel metal2 s 148456 99600 148512 100000 6 instr_write_data[2]
port 117 nsew signal output
rlabel metal2 s 150920 99600 150976 100000 6 instr_write_data[3]
port 118 nsew signal output
rlabel metal2 s 153384 99600 153440 100000 6 instr_write_data[4]
port 119 nsew signal output
rlabel metal2 s 155848 99600 155904 100000 6 instr_write_data[5]
port 120 nsew signal output
rlabel metal2 s 158312 99600 158368 100000 6 instr_write_data[6]
port 121 nsew signal output
rlabel metal2 s 160776 99600 160832 100000 6 instr_write_data[7]
port 122 nsew signal output
rlabel metal2 s 162624 99600 162680 100000 6 instr_write_data[8]
port 123 nsew signal output
rlabel metal2 s 163856 99600 163912 100000 6 instr_write_data[9]
port 124 nsew signal output
rlabel metal2 s 141680 99600 141736 100000 6 instrw_en
port 125 nsew signal output
rlabel metal2 s 144144 99600 144200 100000 6 instrw_en_8bit[0]
port 126 nsew signal output
rlabel metal2 s 146608 99600 146664 100000 6 instrw_en_8bit[1]
port 127 nsew signal output
rlabel metal2 s 149072 99600 149128 100000 6 instrw_en_8bit[2]
port 128 nsew signal output
rlabel metal2 s 151536 99600 151592 100000 6 instrw_en_8bit[3]
port 129 nsew signal output
rlabel metal2 s 154000 99600 154056 100000 6 instrw_en_8bit[4]
port 130 nsew signal output
rlabel metal2 s 156464 99600 156520 100000 6 instrw_en_8bit[5]
port 131 nsew signal output
rlabel metal2 s 158928 99600 158984 100000 6 instrw_en_8bit[6]
port 132 nsew signal output
rlabel metal2 s 161392 99600 161448 100000 6 instrw_en_8bit[7]
port 133 nsew signal output
rlabel metal2 s 6776 99600 6832 100000 6 io_in[0]
port 134 nsew signal input
rlabel metal2 s 25256 99600 25312 100000 6 io_in[10]
port 135 nsew signal input
rlabel metal2 s 27104 99600 27160 100000 6 io_in[11]
port 136 nsew signal input
rlabel metal2 s 28952 99600 29008 100000 6 io_in[12]
port 137 nsew signal input
rlabel metal2 s 30800 99600 30856 100000 6 io_in[13]
port 138 nsew signal input
rlabel metal2 s 32648 99600 32704 100000 6 io_in[14]
port 139 nsew signal input
rlabel metal2 s 34496 99600 34552 100000 6 io_in[15]
port 140 nsew signal input
rlabel metal2 s 36344 99600 36400 100000 6 io_in[16]
port 141 nsew signal input
rlabel metal2 s 38192 99600 38248 100000 6 io_in[17]
port 142 nsew signal input
rlabel metal2 s 40040 99600 40096 100000 6 io_in[18]
port 143 nsew signal input
rlabel metal2 s 41888 99600 41944 100000 6 io_in[19]
port 144 nsew signal input
rlabel metal2 s 8624 99600 8680 100000 6 io_in[1]
port 145 nsew signal input
rlabel metal2 s 43736 99600 43792 100000 6 io_in[20]
port 146 nsew signal input
rlabel metal2 s 45584 99600 45640 100000 6 io_in[21]
port 147 nsew signal input
rlabel metal2 s 47432 99600 47488 100000 6 io_in[22]
port 148 nsew signal input
rlabel metal2 s 49280 99600 49336 100000 6 io_in[23]
port 149 nsew signal input
rlabel metal2 s 51128 99600 51184 100000 6 io_in[24]
port 150 nsew signal input
rlabel metal2 s 52976 99600 53032 100000 6 io_in[25]
port 151 nsew signal input
rlabel metal2 s 54824 99600 54880 100000 6 io_in[26]
port 152 nsew signal input
rlabel metal2 s 56672 99600 56728 100000 6 io_in[27]
port 153 nsew signal input
rlabel metal2 s 58520 99600 58576 100000 6 io_in[28]
port 154 nsew signal input
rlabel metal2 s 60368 99600 60424 100000 6 io_in[29]
port 155 nsew signal input
rlabel metal2 s 10472 99600 10528 100000 6 io_in[2]
port 156 nsew signal input
rlabel metal2 s 62216 99600 62272 100000 6 io_in[30]
port 157 nsew signal input
rlabel metal2 s 64064 99600 64120 100000 6 io_in[31]
port 158 nsew signal input
rlabel metal2 s 65912 99600 65968 100000 6 io_in[32]
port 159 nsew signal input
rlabel metal2 s 67760 99600 67816 100000 6 io_in[33]
port 160 nsew signal input
rlabel metal2 s 69608 99600 69664 100000 6 io_in[34]
port 161 nsew signal input
rlabel metal2 s 71456 99600 71512 100000 6 io_in[35]
port 162 nsew signal input
rlabel metal2 s 73304 99600 73360 100000 6 io_in[36]
port 163 nsew signal input
rlabel metal2 s 75152 99600 75208 100000 6 io_in[37]
port 164 nsew signal input
rlabel metal2 s 12320 99600 12376 100000 6 io_in[3]
port 165 nsew signal input
rlabel metal2 s 14168 99600 14224 100000 6 io_in[4]
port 166 nsew signal input
rlabel metal2 s 16016 99600 16072 100000 6 io_in[5]
port 167 nsew signal input
rlabel metal2 s 17864 99600 17920 100000 6 io_in[6]
port 168 nsew signal input
rlabel metal2 s 19712 99600 19768 100000 6 io_in[7]
port 169 nsew signal input
rlabel metal2 s 21560 99600 21616 100000 6 io_in[8]
port 170 nsew signal input
rlabel metal2 s 23408 99600 23464 100000 6 io_in[9]
port 171 nsew signal input
rlabel metal2 s 7392 99600 7448 100000 6 io_oeb[0]
port 172 nsew signal output
rlabel metal2 s 25872 99600 25928 100000 6 io_oeb[10]
port 173 nsew signal output
rlabel metal2 s 27720 99600 27776 100000 6 io_oeb[11]
port 174 nsew signal output
rlabel metal2 s 29568 99600 29624 100000 6 io_oeb[12]
port 175 nsew signal output
rlabel metal2 s 31416 99600 31472 100000 6 io_oeb[13]
port 176 nsew signal output
rlabel metal2 s 33264 99600 33320 100000 6 io_oeb[14]
port 177 nsew signal output
rlabel metal2 s 35112 99600 35168 100000 6 io_oeb[15]
port 178 nsew signal output
rlabel metal2 s 36960 99600 37016 100000 6 io_oeb[16]
port 179 nsew signal output
rlabel metal2 s 38808 99600 38864 100000 6 io_oeb[17]
port 180 nsew signal output
rlabel metal2 s 40656 99600 40712 100000 6 io_oeb[18]
port 181 nsew signal output
rlabel metal2 s 42504 99600 42560 100000 6 io_oeb[19]
port 182 nsew signal output
rlabel metal2 s 9240 99600 9296 100000 6 io_oeb[1]
port 183 nsew signal output
rlabel metal2 s 44352 99600 44408 100000 6 io_oeb[20]
port 184 nsew signal output
rlabel metal2 s 46200 99600 46256 100000 6 io_oeb[21]
port 185 nsew signal output
rlabel metal2 s 48048 99600 48104 100000 6 io_oeb[22]
port 186 nsew signal output
rlabel metal2 s 49896 99600 49952 100000 6 io_oeb[23]
port 187 nsew signal output
rlabel metal2 s 51744 99600 51800 100000 6 io_oeb[24]
port 188 nsew signal output
rlabel metal2 s 53592 99600 53648 100000 6 io_oeb[25]
port 189 nsew signal output
rlabel metal2 s 55440 99600 55496 100000 6 io_oeb[26]
port 190 nsew signal output
rlabel metal2 s 57288 99600 57344 100000 6 io_oeb[27]
port 191 nsew signal output
rlabel metal2 s 59136 99600 59192 100000 6 io_oeb[28]
port 192 nsew signal output
rlabel metal2 s 60984 99600 61040 100000 6 io_oeb[29]
port 193 nsew signal output
rlabel metal2 s 11088 99600 11144 100000 6 io_oeb[2]
port 194 nsew signal output
rlabel metal2 s 62832 99600 62888 100000 6 io_oeb[30]
port 195 nsew signal output
rlabel metal2 s 64680 99600 64736 100000 6 io_oeb[31]
port 196 nsew signal output
rlabel metal2 s 66528 99600 66584 100000 6 io_oeb[32]
port 197 nsew signal output
rlabel metal2 s 68376 99600 68432 100000 6 io_oeb[33]
port 198 nsew signal output
rlabel metal2 s 70224 99600 70280 100000 6 io_oeb[34]
port 199 nsew signal output
rlabel metal2 s 72072 99600 72128 100000 6 io_oeb[35]
port 200 nsew signal output
rlabel metal2 s 73920 99600 73976 100000 6 io_oeb[36]
port 201 nsew signal output
rlabel metal2 s 75768 99600 75824 100000 6 io_oeb[37]
port 202 nsew signal output
rlabel metal2 s 12936 99600 12992 100000 6 io_oeb[3]
port 203 nsew signal output
rlabel metal2 s 14784 99600 14840 100000 6 io_oeb[4]
port 204 nsew signal output
rlabel metal2 s 16632 99600 16688 100000 6 io_oeb[5]
port 205 nsew signal output
rlabel metal2 s 18480 99600 18536 100000 6 io_oeb[6]
port 206 nsew signal output
rlabel metal2 s 20328 99600 20384 100000 6 io_oeb[7]
port 207 nsew signal output
rlabel metal2 s 22176 99600 22232 100000 6 io_oeb[8]
port 208 nsew signal output
rlabel metal2 s 24024 99600 24080 100000 6 io_oeb[9]
port 209 nsew signal output
rlabel metal2 s 8008 99600 8064 100000 6 io_out[0]
port 210 nsew signal output
rlabel metal2 s 26488 99600 26544 100000 6 io_out[10]
port 211 nsew signal output
rlabel metal2 s 28336 99600 28392 100000 6 io_out[11]
port 212 nsew signal output
rlabel metal2 s 30184 99600 30240 100000 6 io_out[12]
port 213 nsew signal output
rlabel metal2 s 32032 99600 32088 100000 6 io_out[13]
port 214 nsew signal output
rlabel metal2 s 33880 99600 33936 100000 6 io_out[14]
port 215 nsew signal output
rlabel metal2 s 35728 99600 35784 100000 6 io_out[15]
port 216 nsew signal output
rlabel metal2 s 37576 99600 37632 100000 6 io_out[16]
port 217 nsew signal output
rlabel metal2 s 39424 99600 39480 100000 6 io_out[17]
port 218 nsew signal output
rlabel metal2 s 41272 99600 41328 100000 6 io_out[18]
port 219 nsew signal output
rlabel metal2 s 43120 99600 43176 100000 6 io_out[19]
port 220 nsew signal output
rlabel metal2 s 9856 99600 9912 100000 6 io_out[1]
port 221 nsew signal output
rlabel metal2 s 44968 99600 45024 100000 6 io_out[20]
port 222 nsew signal output
rlabel metal2 s 46816 99600 46872 100000 6 io_out[21]
port 223 nsew signal output
rlabel metal2 s 48664 99600 48720 100000 6 io_out[22]
port 224 nsew signal output
rlabel metal2 s 50512 99600 50568 100000 6 io_out[23]
port 225 nsew signal output
rlabel metal2 s 52360 99600 52416 100000 6 io_out[24]
port 226 nsew signal output
rlabel metal2 s 54208 99600 54264 100000 6 io_out[25]
port 227 nsew signal output
rlabel metal2 s 56056 99600 56112 100000 6 io_out[26]
port 228 nsew signal output
rlabel metal2 s 57904 99600 57960 100000 6 io_out[27]
port 229 nsew signal output
rlabel metal2 s 59752 99600 59808 100000 6 io_out[28]
port 230 nsew signal output
rlabel metal2 s 61600 99600 61656 100000 6 io_out[29]
port 231 nsew signal output
rlabel metal2 s 11704 99600 11760 100000 6 io_out[2]
port 232 nsew signal output
rlabel metal2 s 63448 99600 63504 100000 6 io_out[30]
port 233 nsew signal output
rlabel metal2 s 65296 99600 65352 100000 6 io_out[31]
port 234 nsew signal output
rlabel metal2 s 67144 99600 67200 100000 6 io_out[32]
port 235 nsew signal output
rlabel metal2 s 68992 99600 69048 100000 6 io_out[33]
port 236 nsew signal output
rlabel metal2 s 70840 99600 70896 100000 6 io_out[34]
port 237 nsew signal output
rlabel metal2 s 72688 99600 72744 100000 6 io_out[35]
port 238 nsew signal output
rlabel metal2 s 74536 99600 74592 100000 6 io_out[36]
port 239 nsew signal output
rlabel metal2 s 76384 99600 76440 100000 6 io_out[37]
port 240 nsew signal output
rlabel metal2 s 13552 99600 13608 100000 6 io_out[3]
port 241 nsew signal output
rlabel metal2 s 15400 99600 15456 100000 6 io_out[4]
port 242 nsew signal output
rlabel metal2 s 17248 99600 17304 100000 6 io_out[5]
port 243 nsew signal output
rlabel metal2 s 19096 99600 19152 100000 6 io_out[6]
port 244 nsew signal output
rlabel metal2 s 20944 99600 21000 100000 6 io_out[7]
port 245 nsew signal output
rlabel metal2 s 22792 99600 22848 100000 6 io_out[8]
port 246 nsew signal output
rlabel metal2 s 24640 99600 24696 100000 6 io_out[9]
port 247 nsew signal output
rlabel metal2 s 176288 0 176344 400 6 irq[0]
port 248 nsew signal output
rlabel metal2 s 176624 0 176680 400 6 irq[1]
port 249 nsew signal output
rlabel metal2 s 176960 0 177016 400 6 irq[2]
port 250 nsew signal output
rlabel metal2 s 37520 0 37576 400 6 la_data_in[0]
port 251 nsew signal input
rlabel metal2 s 138320 0 138376 400 6 la_data_in[100]
port 252 nsew signal input
rlabel metal2 s 139328 0 139384 400 6 la_data_in[101]
port 253 nsew signal input
rlabel metal2 s 140336 0 140392 400 6 la_data_in[102]
port 254 nsew signal input
rlabel metal2 s 141344 0 141400 400 6 la_data_in[103]
port 255 nsew signal input
rlabel metal2 s 142352 0 142408 400 6 la_data_in[104]
port 256 nsew signal input
rlabel metal2 s 143360 0 143416 400 6 la_data_in[105]
port 257 nsew signal input
rlabel metal2 s 144368 0 144424 400 6 la_data_in[106]
port 258 nsew signal input
rlabel metal2 s 145376 0 145432 400 6 la_data_in[107]
port 259 nsew signal input
rlabel metal2 s 146384 0 146440 400 6 la_data_in[108]
port 260 nsew signal input
rlabel metal2 s 147392 0 147448 400 6 la_data_in[109]
port 261 nsew signal input
rlabel metal2 s 47600 0 47656 400 6 la_data_in[10]
port 262 nsew signal input
rlabel metal2 s 148400 0 148456 400 6 la_data_in[110]
port 263 nsew signal input
rlabel metal2 s 149408 0 149464 400 6 la_data_in[111]
port 264 nsew signal input
rlabel metal2 s 150416 0 150472 400 6 la_data_in[112]
port 265 nsew signal input
rlabel metal2 s 151424 0 151480 400 6 la_data_in[113]
port 266 nsew signal input
rlabel metal2 s 152432 0 152488 400 6 la_data_in[114]
port 267 nsew signal input
rlabel metal2 s 153440 0 153496 400 6 la_data_in[115]
port 268 nsew signal input
rlabel metal2 s 154448 0 154504 400 6 la_data_in[116]
port 269 nsew signal input
rlabel metal2 s 155456 0 155512 400 6 la_data_in[117]
port 270 nsew signal input
rlabel metal2 s 156464 0 156520 400 6 la_data_in[118]
port 271 nsew signal input
rlabel metal2 s 157472 0 157528 400 6 la_data_in[119]
port 272 nsew signal input
rlabel metal2 s 48608 0 48664 400 6 la_data_in[11]
port 273 nsew signal input
rlabel metal2 s 158480 0 158536 400 6 la_data_in[120]
port 274 nsew signal input
rlabel metal2 s 159488 0 159544 400 6 la_data_in[121]
port 275 nsew signal input
rlabel metal2 s 160496 0 160552 400 6 la_data_in[122]
port 276 nsew signal input
rlabel metal2 s 161504 0 161560 400 6 la_data_in[123]
port 277 nsew signal input
rlabel metal2 s 162512 0 162568 400 6 la_data_in[124]
port 278 nsew signal input
rlabel metal2 s 163520 0 163576 400 6 la_data_in[125]
port 279 nsew signal input
rlabel metal2 s 164528 0 164584 400 6 la_data_in[126]
port 280 nsew signal input
rlabel metal2 s 165536 0 165592 400 6 la_data_in[127]
port 281 nsew signal input
rlabel metal2 s 49616 0 49672 400 6 la_data_in[12]
port 282 nsew signal input
rlabel metal2 s 50624 0 50680 400 6 la_data_in[13]
port 283 nsew signal input
rlabel metal2 s 51632 0 51688 400 6 la_data_in[14]
port 284 nsew signal input
rlabel metal2 s 52640 0 52696 400 6 la_data_in[15]
port 285 nsew signal input
rlabel metal2 s 53648 0 53704 400 6 la_data_in[16]
port 286 nsew signal input
rlabel metal2 s 54656 0 54712 400 6 la_data_in[17]
port 287 nsew signal input
rlabel metal2 s 55664 0 55720 400 6 la_data_in[18]
port 288 nsew signal input
rlabel metal2 s 56672 0 56728 400 6 la_data_in[19]
port 289 nsew signal input
rlabel metal2 s 38528 0 38584 400 6 la_data_in[1]
port 290 nsew signal input
rlabel metal2 s 57680 0 57736 400 6 la_data_in[20]
port 291 nsew signal input
rlabel metal2 s 58688 0 58744 400 6 la_data_in[21]
port 292 nsew signal input
rlabel metal2 s 59696 0 59752 400 6 la_data_in[22]
port 293 nsew signal input
rlabel metal2 s 60704 0 60760 400 6 la_data_in[23]
port 294 nsew signal input
rlabel metal2 s 61712 0 61768 400 6 la_data_in[24]
port 295 nsew signal input
rlabel metal2 s 62720 0 62776 400 6 la_data_in[25]
port 296 nsew signal input
rlabel metal2 s 63728 0 63784 400 6 la_data_in[26]
port 297 nsew signal input
rlabel metal2 s 64736 0 64792 400 6 la_data_in[27]
port 298 nsew signal input
rlabel metal2 s 65744 0 65800 400 6 la_data_in[28]
port 299 nsew signal input
rlabel metal2 s 66752 0 66808 400 6 la_data_in[29]
port 300 nsew signal input
rlabel metal2 s 39536 0 39592 400 6 la_data_in[2]
port 301 nsew signal input
rlabel metal2 s 67760 0 67816 400 6 la_data_in[30]
port 302 nsew signal input
rlabel metal2 s 68768 0 68824 400 6 la_data_in[31]
port 303 nsew signal input
rlabel metal2 s 69776 0 69832 400 6 la_data_in[32]
port 304 nsew signal input
rlabel metal2 s 70784 0 70840 400 6 la_data_in[33]
port 305 nsew signal input
rlabel metal2 s 71792 0 71848 400 6 la_data_in[34]
port 306 nsew signal input
rlabel metal2 s 72800 0 72856 400 6 la_data_in[35]
port 307 nsew signal input
rlabel metal2 s 73808 0 73864 400 6 la_data_in[36]
port 308 nsew signal input
rlabel metal2 s 74816 0 74872 400 6 la_data_in[37]
port 309 nsew signal input
rlabel metal2 s 75824 0 75880 400 6 la_data_in[38]
port 310 nsew signal input
rlabel metal2 s 76832 0 76888 400 6 la_data_in[39]
port 311 nsew signal input
rlabel metal2 s 40544 0 40600 400 6 la_data_in[3]
port 312 nsew signal input
rlabel metal2 s 77840 0 77896 400 6 la_data_in[40]
port 313 nsew signal input
rlabel metal2 s 78848 0 78904 400 6 la_data_in[41]
port 314 nsew signal input
rlabel metal2 s 79856 0 79912 400 6 la_data_in[42]
port 315 nsew signal input
rlabel metal2 s 80864 0 80920 400 6 la_data_in[43]
port 316 nsew signal input
rlabel metal2 s 81872 0 81928 400 6 la_data_in[44]
port 317 nsew signal input
rlabel metal2 s 82880 0 82936 400 6 la_data_in[45]
port 318 nsew signal input
rlabel metal2 s 83888 0 83944 400 6 la_data_in[46]
port 319 nsew signal input
rlabel metal2 s 84896 0 84952 400 6 la_data_in[47]
port 320 nsew signal input
rlabel metal2 s 85904 0 85960 400 6 la_data_in[48]
port 321 nsew signal input
rlabel metal2 s 86912 0 86968 400 6 la_data_in[49]
port 322 nsew signal input
rlabel metal2 s 41552 0 41608 400 6 la_data_in[4]
port 323 nsew signal input
rlabel metal2 s 87920 0 87976 400 6 la_data_in[50]
port 324 nsew signal input
rlabel metal2 s 88928 0 88984 400 6 la_data_in[51]
port 325 nsew signal input
rlabel metal2 s 89936 0 89992 400 6 la_data_in[52]
port 326 nsew signal input
rlabel metal2 s 90944 0 91000 400 6 la_data_in[53]
port 327 nsew signal input
rlabel metal2 s 91952 0 92008 400 6 la_data_in[54]
port 328 nsew signal input
rlabel metal2 s 92960 0 93016 400 6 la_data_in[55]
port 329 nsew signal input
rlabel metal2 s 93968 0 94024 400 6 la_data_in[56]
port 330 nsew signal input
rlabel metal2 s 94976 0 95032 400 6 la_data_in[57]
port 331 nsew signal input
rlabel metal2 s 95984 0 96040 400 6 la_data_in[58]
port 332 nsew signal input
rlabel metal2 s 96992 0 97048 400 6 la_data_in[59]
port 333 nsew signal input
rlabel metal2 s 42560 0 42616 400 6 la_data_in[5]
port 334 nsew signal input
rlabel metal2 s 98000 0 98056 400 6 la_data_in[60]
port 335 nsew signal input
rlabel metal2 s 99008 0 99064 400 6 la_data_in[61]
port 336 nsew signal input
rlabel metal2 s 100016 0 100072 400 6 la_data_in[62]
port 337 nsew signal input
rlabel metal2 s 101024 0 101080 400 6 la_data_in[63]
port 338 nsew signal input
rlabel metal2 s 102032 0 102088 400 6 la_data_in[64]
port 339 nsew signal input
rlabel metal2 s 103040 0 103096 400 6 la_data_in[65]
port 340 nsew signal input
rlabel metal2 s 104048 0 104104 400 6 la_data_in[66]
port 341 nsew signal input
rlabel metal2 s 105056 0 105112 400 6 la_data_in[67]
port 342 nsew signal input
rlabel metal2 s 106064 0 106120 400 6 la_data_in[68]
port 343 nsew signal input
rlabel metal2 s 107072 0 107128 400 6 la_data_in[69]
port 344 nsew signal input
rlabel metal2 s 43568 0 43624 400 6 la_data_in[6]
port 345 nsew signal input
rlabel metal2 s 108080 0 108136 400 6 la_data_in[70]
port 346 nsew signal input
rlabel metal2 s 109088 0 109144 400 6 la_data_in[71]
port 347 nsew signal input
rlabel metal2 s 110096 0 110152 400 6 la_data_in[72]
port 348 nsew signal input
rlabel metal2 s 111104 0 111160 400 6 la_data_in[73]
port 349 nsew signal input
rlabel metal2 s 112112 0 112168 400 6 la_data_in[74]
port 350 nsew signal input
rlabel metal2 s 113120 0 113176 400 6 la_data_in[75]
port 351 nsew signal input
rlabel metal2 s 114128 0 114184 400 6 la_data_in[76]
port 352 nsew signal input
rlabel metal2 s 115136 0 115192 400 6 la_data_in[77]
port 353 nsew signal input
rlabel metal2 s 116144 0 116200 400 6 la_data_in[78]
port 354 nsew signal input
rlabel metal2 s 117152 0 117208 400 6 la_data_in[79]
port 355 nsew signal input
rlabel metal2 s 44576 0 44632 400 6 la_data_in[7]
port 356 nsew signal input
rlabel metal2 s 118160 0 118216 400 6 la_data_in[80]
port 357 nsew signal input
rlabel metal2 s 119168 0 119224 400 6 la_data_in[81]
port 358 nsew signal input
rlabel metal2 s 120176 0 120232 400 6 la_data_in[82]
port 359 nsew signal input
rlabel metal2 s 121184 0 121240 400 6 la_data_in[83]
port 360 nsew signal input
rlabel metal2 s 122192 0 122248 400 6 la_data_in[84]
port 361 nsew signal input
rlabel metal2 s 123200 0 123256 400 6 la_data_in[85]
port 362 nsew signal input
rlabel metal2 s 124208 0 124264 400 6 la_data_in[86]
port 363 nsew signal input
rlabel metal2 s 125216 0 125272 400 6 la_data_in[87]
port 364 nsew signal input
rlabel metal2 s 126224 0 126280 400 6 la_data_in[88]
port 365 nsew signal input
rlabel metal2 s 127232 0 127288 400 6 la_data_in[89]
port 366 nsew signal input
rlabel metal2 s 45584 0 45640 400 6 la_data_in[8]
port 367 nsew signal input
rlabel metal2 s 128240 0 128296 400 6 la_data_in[90]
port 368 nsew signal input
rlabel metal2 s 129248 0 129304 400 6 la_data_in[91]
port 369 nsew signal input
rlabel metal2 s 130256 0 130312 400 6 la_data_in[92]
port 370 nsew signal input
rlabel metal2 s 131264 0 131320 400 6 la_data_in[93]
port 371 nsew signal input
rlabel metal2 s 132272 0 132328 400 6 la_data_in[94]
port 372 nsew signal input
rlabel metal2 s 133280 0 133336 400 6 la_data_in[95]
port 373 nsew signal input
rlabel metal2 s 134288 0 134344 400 6 la_data_in[96]
port 374 nsew signal input
rlabel metal2 s 135296 0 135352 400 6 la_data_in[97]
port 375 nsew signal input
rlabel metal2 s 136304 0 136360 400 6 la_data_in[98]
port 376 nsew signal input
rlabel metal2 s 137312 0 137368 400 6 la_data_in[99]
port 377 nsew signal input
rlabel metal2 s 46592 0 46648 400 6 la_data_in[9]
port 378 nsew signal input
rlabel metal2 s 37856 0 37912 400 6 la_data_out[0]
port 379 nsew signal output
rlabel metal2 s 138656 0 138712 400 6 la_data_out[100]
port 380 nsew signal output
rlabel metal2 s 139664 0 139720 400 6 la_data_out[101]
port 381 nsew signal output
rlabel metal2 s 140672 0 140728 400 6 la_data_out[102]
port 382 nsew signal output
rlabel metal2 s 141680 0 141736 400 6 la_data_out[103]
port 383 nsew signal output
rlabel metal2 s 142688 0 142744 400 6 la_data_out[104]
port 384 nsew signal output
rlabel metal2 s 143696 0 143752 400 6 la_data_out[105]
port 385 nsew signal output
rlabel metal2 s 144704 0 144760 400 6 la_data_out[106]
port 386 nsew signal output
rlabel metal2 s 145712 0 145768 400 6 la_data_out[107]
port 387 nsew signal output
rlabel metal2 s 146720 0 146776 400 6 la_data_out[108]
port 388 nsew signal output
rlabel metal2 s 147728 0 147784 400 6 la_data_out[109]
port 389 nsew signal output
rlabel metal2 s 47936 0 47992 400 6 la_data_out[10]
port 390 nsew signal output
rlabel metal2 s 148736 0 148792 400 6 la_data_out[110]
port 391 nsew signal output
rlabel metal2 s 149744 0 149800 400 6 la_data_out[111]
port 392 nsew signal output
rlabel metal2 s 150752 0 150808 400 6 la_data_out[112]
port 393 nsew signal output
rlabel metal2 s 151760 0 151816 400 6 la_data_out[113]
port 394 nsew signal output
rlabel metal2 s 152768 0 152824 400 6 la_data_out[114]
port 395 nsew signal output
rlabel metal2 s 153776 0 153832 400 6 la_data_out[115]
port 396 nsew signal output
rlabel metal2 s 154784 0 154840 400 6 la_data_out[116]
port 397 nsew signal output
rlabel metal2 s 155792 0 155848 400 6 la_data_out[117]
port 398 nsew signal output
rlabel metal2 s 156800 0 156856 400 6 la_data_out[118]
port 399 nsew signal output
rlabel metal2 s 157808 0 157864 400 6 la_data_out[119]
port 400 nsew signal output
rlabel metal2 s 48944 0 49000 400 6 la_data_out[11]
port 401 nsew signal output
rlabel metal2 s 158816 0 158872 400 6 la_data_out[120]
port 402 nsew signal output
rlabel metal2 s 159824 0 159880 400 6 la_data_out[121]
port 403 nsew signal output
rlabel metal2 s 160832 0 160888 400 6 la_data_out[122]
port 404 nsew signal output
rlabel metal2 s 161840 0 161896 400 6 la_data_out[123]
port 405 nsew signal output
rlabel metal2 s 162848 0 162904 400 6 la_data_out[124]
port 406 nsew signal output
rlabel metal2 s 163856 0 163912 400 6 la_data_out[125]
port 407 nsew signal output
rlabel metal2 s 164864 0 164920 400 6 la_data_out[126]
port 408 nsew signal output
rlabel metal2 s 165872 0 165928 400 6 la_data_out[127]
port 409 nsew signal output
rlabel metal2 s 49952 0 50008 400 6 la_data_out[12]
port 410 nsew signal output
rlabel metal2 s 50960 0 51016 400 6 la_data_out[13]
port 411 nsew signal output
rlabel metal2 s 51968 0 52024 400 6 la_data_out[14]
port 412 nsew signal output
rlabel metal2 s 52976 0 53032 400 6 la_data_out[15]
port 413 nsew signal output
rlabel metal2 s 53984 0 54040 400 6 la_data_out[16]
port 414 nsew signal output
rlabel metal2 s 54992 0 55048 400 6 la_data_out[17]
port 415 nsew signal output
rlabel metal2 s 56000 0 56056 400 6 la_data_out[18]
port 416 nsew signal output
rlabel metal2 s 57008 0 57064 400 6 la_data_out[19]
port 417 nsew signal output
rlabel metal2 s 38864 0 38920 400 6 la_data_out[1]
port 418 nsew signal output
rlabel metal2 s 58016 0 58072 400 6 la_data_out[20]
port 419 nsew signal output
rlabel metal2 s 59024 0 59080 400 6 la_data_out[21]
port 420 nsew signal output
rlabel metal2 s 60032 0 60088 400 6 la_data_out[22]
port 421 nsew signal output
rlabel metal2 s 61040 0 61096 400 6 la_data_out[23]
port 422 nsew signal output
rlabel metal2 s 62048 0 62104 400 6 la_data_out[24]
port 423 nsew signal output
rlabel metal2 s 63056 0 63112 400 6 la_data_out[25]
port 424 nsew signal output
rlabel metal2 s 64064 0 64120 400 6 la_data_out[26]
port 425 nsew signal output
rlabel metal2 s 65072 0 65128 400 6 la_data_out[27]
port 426 nsew signal output
rlabel metal2 s 66080 0 66136 400 6 la_data_out[28]
port 427 nsew signal output
rlabel metal2 s 67088 0 67144 400 6 la_data_out[29]
port 428 nsew signal output
rlabel metal2 s 39872 0 39928 400 6 la_data_out[2]
port 429 nsew signal output
rlabel metal2 s 68096 0 68152 400 6 la_data_out[30]
port 430 nsew signal output
rlabel metal2 s 69104 0 69160 400 6 la_data_out[31]
port 431 nsew signal output
rlabel metal2 s 70112 0 70168 400 6 la_data_out[32]
port 432 nsew signal output
rlabel metal2 s 71120 0 71176 400 6 la_data_out[33]
port 433 nsew signal output
rlabel metal2 s 72128 0 72184 400 6 la_data_out[34]
port 434 nsew signal output
rlabel metal2 s 73136 0 73192 400 6 la_data_out[35]
port 435 nsew signal output
rlabel metal2 s 74144 0 74200 400 6 la_data_out[36]
port 436 nsew signal output
rlabel metal2 s 75152 0 75208 400 6 la_data_out[37]
port 437 nsew signal output
rlabel metal2 s 76160 0 76216 400 6 la_data_out[38]
port 438 nsew signal output
rlabel metal2 s 77168 0 77224 400 6 la_data_out[39]
port 439 nsew signal output
rlabel metal2 s 40880 0 40936 400 6 la_data_out[3]
port 440 nsew signal output
rlabel metal2 s 78176 0 78232 400 6 la_data_out[40]
port 441 nsew signal output
rlabel metal2 s 79184 0 79240 400 6 la_data_out[41]
port 442 nsew signal output
rlabel metal2 s 80192 0 80248 400 6 la_data_out[42]
port 443 nsew signal output
rlabel metal2 s 81200 0 81256 400 6 la_data_out[43]
port 444 nsew signal output
rlabel metal2 s 82208 0 82264 400 6 la_data_out[44]
port 445 nsew signal output
rlabel metal2 s 83216 0 83272 400 6 la_data_out[45]
port 446 nsew signal output
rlabel metal2 s 84224 0 84280 400 6 la_data_out[46]
port 447 nsew signal output
rlabel metal2 s 85232 0 85288 400 6 la_data_out[47]
port 448 nsew signal output
rlabel metal2 s 86240 0 86296 400 6 la_data_out[48]
port 449 nsew signal output
rlabel metal2 s 87248 0 87304 400 6 la_data_out[49]
port 450 nsew signal output
rlabel metal2 s 41888 0 41944 400 6 la_data_out[4]
port 451 nsew signal output
rlabel metal2 s 88256 0 88312 400 6 la_data_out[50]
port 452 nsew signal output
rlabel metal2 s 89264 0 89320 400 6 la_data_out[51]
port 453 nsew signal output
rlabel metal2 s 90272 0 90328 400 6 la_data_out[52]
port 454 nsew signal output
rlabel metal2 s 91280 0 91336 400 6 la_data_out[53]
port 455 nsew signal output
rlabel metal2 s 92288 0 92344 400 6 la_data_out[54]
port 456 nsew signal output
rlabel metal2 s 93296 0 93352 400 6 la_data_out[55]
port 457 nsew signal output
rlabel metal2 s 94304 0 94360 400 6 la_data_out[56]
port 458 nsew signal output
rlabel metal2 s 95312 0 95368 400 6 la_data_out[57]
port 459 nsew signal output
rlabel metal2 s 96320 0 96376 400 6 la_data_out[58]
port 460 nsew signal output
rlabel metal2 s 97328 0 97384 400 6 la_data_out[59]
port 461 nsew signal output
rlabel metal2 s 42896 0 42952 400 6 la_data_out[5]
port 462 nsew signal output
rlabel metal2 s 98336 0 98392 400 6 la_data_out[60]
port 463 nsew signal output
rlabel metal2 s 99344 0 99400 400 6 la_data_out[61]
port 464 nsew signal output
rlabel metal2 s 100352 0 100408 400 6 la_data_out[62]
port 465 nsew signal output
rlabel metal2 s 101360 0 101416 400 6 la_data_out[63]
port 466 nsew signal output
rlabel metal2 s 102368 0 102424 400 6 la_data_out[64]
port 467 nsew signal output
rlabel metal2 s 103376 0 103432 400 6 la_data_out[65]
port 468 nsew signal output
rlabel metal2 s 104384 0 104440 400 6 la_data_out[66]
port 469 nsew signal output
rlabel metal2 s 105392 0 105448 400 6 la_data_out[67]
port 470 nsew signal output
rlabel metal2 s 106400 0 106456 400 6 la_data_out[68]
port 471 nsew signal output
rlabel metal2 s 107408 0 107464 400 6 la_data_out[69]
port 472 nsew signal output
rlabel metal2 s 43904 0 43960 400 6 la_data_out[6]
port 473 nsew signal output
rlabel metal2 s 108416 0 108472 400 6 la_data_out[70]
port 474 nsew signal output
rlabel metal2 s 109424 0 109480 400 6 la_data_out[71]
port 475 nsew signal output
rlabel metal2 s 110432 0 110488 400 6 la_data_out[72]
port 476 nsew signal output
rlabel metal2 s 111440 0 111496 400 6 la_data_out[73]
port 477 nsew signal output
rlabel metal2 s 112448 0 112504 400 6 la_data_out[74]
port 478 nsew signal output
rlabel metal2 s 113456 0 113512 400 6 la_data_out[75]
port 479 nsew signal output
rlabel metal2 s 114464 0 114520 400 6 la_data_out[76]
port 480 nsew signal output
rlabel metal2 s 115472 0 115528 400 6 la_data_out[77]
port 481 nsew signal output
rlabel metal2 s 116480 0 116536 400 6 la_data_out[78]
port 482 nsew signal output
rlabel metal2 s 117488 0 117544 400 6 la_data_out[79]
port 483 nsew signal output
rlabel metal2 s 44912 0 44968 400 6 la_data_out[7]
port 484 nsew signal output
rlabel metal2 s 118496 0 118552 400 6 la_data_out[80]
port 485 nsew signal output
rlabel metal2 s 119504 0 119560 400 6 la_data_out[81]
port 486 nsew signal output
rlabel metal2 s 120512 0 120568 400 6 la_data_out[82]
port 487 nsew signal output
rlabel metal2 s 121520 0 121576 400 6 la_data_out[83]
port 488 nsew signal output
rlabel metal2 s 122528 0 122584 400 6 la_data_out[84]
port 489 nsew signal output
rlabel metal2 s 123536 0 123592 400 6 la_data_out[85]
port 490 nsew signal output
rlabel metal2 s 124544 0 124600 400 6 la_data_out[86]
port 491 nsew signal output
rlabel metal2 s 125552 0 125608 400 6 la_data_out[87]
port 492 nsew signal output
rlabel metal2 s 126560 0 126616 400 6 la_data_out[88]
port 493 nsew signal output
rlabel metal2 s 127568 0 127624 400 6 la_data_out[89]
port 494 nsew signal output
rlabel metal2 s 45920 0 45976 400 6 la_data_out[8]
port 495 nsew signal output
rlabel metal2 s 128576 0 128632 400 6 la_data_out[90]
port 496 nsew signal output
rlabel metal2 s 129584 0 129640 400 6 la_data_out[91]
port 497 nsew signal output
rlabel metal2 s 130592 0 130648 400 6 la_data_out[92]
port 498 nsew signal output
rlabel metal2 s 131600 0 131656 400 6 la_data_out[93]
port 499 nsew signal output
rlabel metal2 s 132608 0 132664 400 6 la_data_out[94]
port 500 nsew signal output
rlabel metal2 s 133616 0 133672 400 6 la_data_out[95]
port 501 nsew signal output
rlabel metal2 s 134624 0 134680 400 6 la_data_out[96]
port 502 nsew signal output
rlabel metal2 s 135632 0 135688 400 6 la_data_out[97]
port 503 nsew signal output
rlabel metal2 s 136640 0 136696 400 6 la_data_out[98]
port 504 nsew signal output
rlabel metal2 s 137648 0 137704 400 6 la_data_out[99]
port 505 nsew signal output
rlabel metal2 s 46928 0 46984 400 6 la_data_out[9]
port 506 nsew signal output
rlabel metal2 s 38192 0 38248 400 6 la_oenb[0]
port 507 nsew signal input
rlabel metal2 s 138992 0 139048 400 6 la_oenb[100]
port 508 nsew signal input
rlabel metal2 s 140000 0 140056 400 6 la_oenb[101]
port 509 nsew signal input
rlabel metal2 s 141008 0 141064 400 6 la_oenb[102]
port 510 nsew signal input
rlabel metal2 s 142016 0 142072 400 6 la_oenb[103]
port 511 nsew signal input
rlabel metal2 s 143024 0 143080 400 6 la_oenb[104]
port 512 nsew signal input
rlabel metal2 s 144032 0 144088 400 6 la_oenb[105]
port 513 nsew signal input
rlabel metal2 s 145040 0 145096 400 6 la_oenb[106]
port 514 nsew signal input
rlabel metal2 s 146048 0 146104 400 6 la_oenb[107]
port 515 nsew signal input
rlabel metal2 s 147056 0 147112 400 6 la_oenb[108]
port 516 nsew signal input
rlabel metal2 s 148064 0 148120 400 6 la_oenb[109]
port 517 nsew signal input
rlabel metal2 s 48272 0 48328 400 6 la_oenb[10]
port 518 nsew signal input
rlabel metal2 s 149072 0 149128 400 6 la_oenb[110]
port 519 nsew signal input
rlabel metal2 s 150080 0 150136 400 6 la_oenb[111]
port 520 nsew signal input
rlabel metal2 s 151088 0 151144 400 6 la_oenb[112]
port 521 nsew signal input
rlabel metal2 s 152096 0 152152 400 6 la_oenb[113]
port 522 nsew signal input
rlabel metal2 s 153104 0 153160 400 6 la_oenb[114]
port 523 nsew signal input
rlabel metal2 s 154112 0 154168 400 6 la_oenb[115]
port 524 nsew signal input
rlabel metal2 s 155120 0 155176 400 6 la_oenb[116]
port 525 nsew signal input
rlabel metal2 s 156128 0 156184 400 6 la_oenb[117]
port 526 nsew signal input
rlabel metal2 s 157136 0 157192 400 6 la_oenb[118]
port 527 nsew signal input
rlabel metal2 s 158144 0 158200 400 6 la_oenb[119]
port 528 nsew signal input
rlabel metal2 s 49280 0 49336 400 6 la_oenb[11]
port 529 nsew signal input
rlabel metal2 s 159152 0 159208 400 6 la_oenb[120]
port 530 nsew signal input
rlabel metal2 s 160160 0 160216 400 6 la_oenb[121]
port 531 nsew signal input
rlabel metal2 s 161168 0 161224 400 6 la_oenb[122]
port 532 nsew signal input
rlabel metal2 s 162176 0 162232 400 6 la_oenb[123]
port 533 nsew signal input
rlabel metal2 s 163184 0 163240 400 6 la_oenb[124]
port 534 nsew signal input
rlabel metal2 s 164192 0 164248 400 6 la_oenb[125]
port 535 nsew signal input
rlabel metal2 s 165200 0 165256 400 6 la_oenb[126]
port 536 nsew signal input
rlabel metal2 s 166208 0 166264 400 6 la_oenb[127]
port 537 nsew signal input
rlabel metal2 s 50288 0 50344 400 6 la_oenb[12]
port 538 nsew signal input
rlabel metal2 s 51296 0 51352 400 6 la_oenb[13]
port 539 nsew signal input
rlabel metal2 s 52304 0 52360 400 6 la_oenb[14]
port 540 nsew signal input
rlabel metal2 s 53312 0 53368 400 6 la_oenb[15]
port 541 nsew signal input
rlabel metal2 s 54320 0 54376 400 6 la_oenb[16]
port 542 nsew signal input
rlabel metal2 s 55328 0 55384 400 6 la_oenb[17]
port 543 nsew signal input
rlabel metal2 s 56336 0 56392 400 6 la_oenb[18]
port 544 nsew signal input
rlabel metal2 s 57344 0 57400 400 6 la_oenb[19]
port 545 nsew signal input
rlabel metal2 s 39200 0 39256 400 6 la_oenb[1]
port 546 nsew signal input
rlabel metal2 s 58352 0 58408 400 6 la_oenb[20]
port 547 nsew signal input
rlabel metal2 s 59360 0 59416 400 6 la_oenb[21]
port 548 nsew signal input
rlabel metal2 s 60368 0 60424 400 6 la_oenb[22]
port 549 nsew signal input
rlabel metal2 s 61376 0 61432 400 6 la_oenb[23]
port 550 nsew signal input
rlabel metal2 s 62384 0 62440 400 6 la_oenb[24]
port 551 nsew signal input
rlabel metal2 s 63392 0 63448 400 6 la_oenb[25]
port 552 nsew signal input
rlabel metal2 s 64400 0 64456 400 6 la_oenb[26]
port 553 nsew signal input
rlabel metal2 s 65408 0 65464 400 6 la_oenb[27]
port 554 nsew signal input
rlabel metal2 s 66416 0 66472 400 6 la_oenb[28]
port 555 nsew signal input
rlabel metal2 s 67424 0 67480 400 6 la_oenb[29]
port 556 nsew signal input
rlabel metal2 s 40208 0 40264 400 6 la_oenb[2]
port 557 nsew signal input
rlabel metal2 s 68432 0 68488 400 6 la_oenb[30]
port 558 nsew signal input
rlabel metal2 s 69440 0 69496 400 6 la_oenb[31]
port 559 nsew signal input
rlabel metal2 s 70448 0 70504 400 6 la_oenb[32]
port 560 nsew signal input
rlabel metal2 s 71456 0 71512 400 6 la_oenb[33]
port 561 nsew signal input
rlabel metal2 s 72464 0 72520 400 6 la_oenb[34]
port 562 nsew signal input
rlabel metal2 s 73472 0 73528 400 6 la_oenb[35]
port 563 nsew signal input
rlabel metal2 s 74480 0 74536 400 6 la_oenb[36]
port 564 nsew signal input
rlabel metal2 s 75488 0 75544 400 6 la_oenb[37]
port 565 nsew signal input
rlabel metal2 s 76496 0 76552 400 6 la_oenb[38]
port 566 nsew signal input
rlabel metal2 s 77504 0 77560 400 6 la_oenb[39]
port 567 nsew signal input
rlabel metal2 s 41216 0 41272 400 6 la_oenb[3]
port 568 nsew signal input
rlabel metal2 s 78512 0 78568 400 6 la_oenb[40]
port 569 nsew signal input
rlabel metal2 s 79520 0 79576 400 6 la_oenb[41]
port 570 nsew signal input
rlabel metal2 s 80528 0 80584 400 6 la_oenb[42]
port 571 nsew signal input
rlabel metal2 s 81536 0 81592 400 6 la_oenb[43]
port 572 nsew signal input
rlabel metal2 s 82544 0 82600 400 6 la_oenb[44]
port 573 nsew signal input
rlabel metal2 s 83552 0 83608 400 6 la_oenb[45]
port 574 nsew signal input
rlabel metal2 s 84560 0 84616 400 6 la_oenb[46]
port 575 nsew signal input
rlabel metal2 s 85568 0 85624 400 6 la_oenb[47]
port 576 nsew signal input
rlabel metal2 s 86576 0 86632 400 6 la_oenb[48]
port 577 nsew signal input
rlabel metal2 s 87584 0 87640 400 6 la_oenb[49]
port 578 nsew signal input
rlabel metal2 s 42224 0 42280 400 6 la_oenb[4]
port 579 nsew signal input
rlabel metal2 s 88592 0 88648 400 6 la_oenb[50]
port 580 nsew signal input
rlabel metal2 s 89600 0 89656 400 6 la_oenb[51]
port 581 nsew signal input
rlabel metal2 s 90608 0 90664 400 6 la_oenb[52]
port 582 nsew signal input
rlabel metal2 s 91616 0 91672 400 6 la_oenb[53]
port 583 nsew signal input
rlabel metal2 s 92624 0 92680 400 6 la_oenb[54]
port 584 nsew signal input
rlabel metal2 s 93632 0 93688 400 6 la_oenb[55]
port 585 nsew signal input
rlabel metal2 s 94640 0 94696 400 6 la_oenb[56]
port 586 nsew signal input
rlabel metal2 s 95648 0 95704 400 6 la_oenb[57]
port 587 nsew signal input
rlabel metal2 s 96656 0 96712 400 6 la_oenb[58]
port 588 nsew signal input
rlabel metal2 s 97664 0 97720 400 6 la_oenb[59]
port 589 nsew signal input
rlabel metal2 s 43232 0 43288 400 6 la_oenb[5]
port 590 nsew signal input
rlabel metal2 s 98672 0 98728 400 6 la_oenb[60]
port 591 nsew signal input
rlabel metal2 s 99680 0 99736 400 6 la_oenb[61]
port 592 nsew signal input
rlabel metal2 s 100688 0 100744 400 6 la_oenb[62]
port 593 nsew signal input
rlabel metal2 s 101696 0 101752 400 6 la_oenb[63]
port 594 nsew signal input
rlabel metal2 s 102704 0 102760 400 6 la_oenb[64]
port 595 nsew signal input
rlabel metal2 s 103712 0 103768 400 6 la_oenb[65]
port 596 nsew signal input
rlabel metal2 s 104720 0 104776 400 6 la_oenb[66]
port 597 nsew signal input
rlabel metal2 s 105728 0 105784 400 6 la_oenb[67]
port 598 nsew signal input
rlabel metal2 s 106736 0 106792 400 6 la_oenb[68]
port 599 nsew signal input
rlabel metal2 s 107744 0 107800 400 6 la_oenb[69]
port 600 nsew signal input
rlabel metal2 s 44240 0 44296 400 6 la_oenb[6]
port 601 nsew signal input
rlabel metal2 s 108752 0 108808 400 6 la_oenb[70]
port 602 nsew signal input
rlabel metal2 s 109760 0 109816 400 6 la_oenb[71]
port 603 nsew signal input
rlabel metal2 s 110768 0 110824 400 6 la_oenb[72]
port 604 nsew signal input
rlabel metal2 s 111776 0 111832 400 6 la_oenb[73]
port 605 nsew signal input
rlabel metal2 s 112784 0 112840 400 6 la_oenb[74]
port 606 nsew signal input
rlabel metal2 s 113792 0 113848 400 6 la_oenb[75]
port 607 nsew signal input
rlabel metal2 s 114800 0 114856 400 6 la_oenb[76]
port 608 nsew signal input
rlabel metal2 s 115808 0 115864 400 6 la_oenb[77]
port 609 nsew signal input
rlabel metal2 s 116816 0 116872 400 6 la_oenb[78]
port 610 nsew signal input
rlabel metal2 s 117824 0 117880 400 6 la_oenb[79]
port 611 nsew signal input
rlabel metal2 s 45248 0 45304 400 6 la_oenb[7]
port 612 nsew signal input
rlabel metal2 s 118832 0 118888 400 6 la_oenb[80]
port 613 nsew signal input
rlabel metal2 s 119840 0 119896 400 6 la_oenb[81]
port 614 nsew signal input
rlabel metal2 s 120848 0 120904 400 6 la_oenb[82]
port 615 nsew signal input
rlabel metal2 s 121856 0 121912 400 6 la_oenb[83]
port 616 nsew signal input
rlabel metal2 s 122864 0 122920 400 6 la_oenb[84]
port 617 nsew signal input
rlabel metal2 s 123872 0 123928 400 6 la_oenb[85]
port 618 nsew signal input
rlabel metal2 s 124880 0 124936 400 6 la_oenb[86]
port 619 nsew signal input
rlabel metal2 s 125888 0 125944 400 6 la_oenb[87]
port 620 nsew signal input
rlabel metal2 s 126896 0 126952 400 6 la_oenb[88]
port 621 nsew signal input
rlabel metal2 s 127904 0 127960 400 6 la_oenb[89]
port 622 nsew signal input
rlabel metal2 s 46256 0 46312 400 6 la_oenb[8]
port 623 nsew signal input
rlabel metal2 s 128912 0 128968 400 6 la_oenb[90]
port 624 nsew signal input
rlabel metal2 s 129920 0 129976 400 6 la_oenb[91]
port 625 nsew signal input
rlabel metal2 s 130928 0 130984 400 6 la_oenb[92]
port 626 nsew signal input
rlabel metal2 s 131936 0 131992 400 6 la_oenb[93]
port 627 nsew signal input
rlabel metal2 s 132944 0 133000 400 6 la_oenb[94]
port 628 nsew signal input
rlabel metal2 s 133952 0 134008 400 6 la_oenb[95]
port 629 nsew signal input
rlabel metal2 s 134960 0 135016 400 6 la_oenb[96]
port 630 nsew signal input
rlabel metal2 s 135968 0 136024 400 6 la_oenb[97]
port 631 nsew signal input
rlabel metal2 s 136976 0 137032 400 6 la_oenb[98]
port 632 nsew signal input
rlabel metal2 s 137984 0 138040 400 6 la_oenb[99]
port 633 nsew signal input
rlabel metal2 s 47264 0 47320 400 6 la_oenb[9]
port 634 nsew signal input
rlabel metal2 s 177968 0 178024 400 6 reset
port 635 nsew signal output
rlabel metal2 s 177632 0 177688 400 6 start
port 636 nsew signal output
rlabel metal2 s 77616 99600 77672 100000 6 uP_data_mem_addr[0]
port 637 nsew signal input
rlabel metal2 s 80080 99600 80136 100000 6 uP_data_mem_addr[1]
port 638 nsew signal input
rlabel metal2 s 82544 99600 82600 100000 6 uP_data_mem_addr[2]
port 639 nsew signal input
rlabel metal2 s 85008 99600 85064 100000 6 uP_data_mem_addr[3]
port 640 nsew signal input
rlabel metal2 s 87472 99600 87528 100000 6 uP_data_mem_addr[4]
port 641 nsew signal input
rlabel metal2 s 89936 99600 89992 100000 6 uP_data_mem_addr[5]
port 642 nsew signal input
rlabel metal2 s 92400 99600 92456 100000 6 uP_data_mem_addr[6]
port 643 nsew signal input
rlabel metal2 s 94864 99600 94920 100000 6 uP_data_mem_addr[7]
port 644 nsew signal input
rlabel metal2 s 77000 99600 77056 100000 6 uP_dataw_en
port 645 nsew signal input
rlabel metal2 s 78232 99600 78288 100000 6 uP_instr[0]
port 646 nsew signal output
rlabel metal2 s 101024 99600 101080 100000 6 uP_instr[10]
port 647 nsew signal output
rlabel metal2 s 102872 99600 102928 100000 6 uP_instr[11]
port 648 nsew signal output
rlabel metal2 s 104720 99600 104776 100000 6 uP_instr[12]
port 649 nsew signal output
rlabel metal2 s 106568 99600 106624 100000 6 uP_instr[13]
port 650 nsew signal output
rlabel metal2 s 107800 99600 107856 100000 6 uP_instr[14]
port 651 nsew signal output
rlabel metal2 s 109032 99600 109088 100000 6 uP_instr[15]
port 652 nsew signal output
rlabel metal2 s 80696 99600 80752 100000 6 uP_instr[1]
port 653 nsew signal output
rlabel metal2 s 83160 99600 83216 100000 6 uP_instr[2]
port 654 nsew signal output
rlabel metal2 s 85624 99600 85680 100000 6 uP_instr[3]
port 655 nsew signal output
rlabel metal2 s 88088 99600 88144 100000 6 uP_instr[4]
port 656 nsew signal output
rlabel metal2 s 90552 99600 90608 100000 6 uP_instr[5]
port 657 nsew signal output
rlabel metal2 s 93016 99600 93072 100000 6 uP_instr[6]
port 658 nsew signal output
rlabel metal2 s 95480 99600 95536 100000 6 uP_instr[7]
port 659 nsew signal output
rlabel metal2 s 97328 99600 97384 100000 6 uP_instr[8]
port 660 nsew signal output
rlabel metal2 s 99176 99600 99232 100000 6 uP_instr[9]
port 661 nsew signal output
rlabel metal2 s 78848 99600 78904 100000 6 uP_instr_mem_addr[0]
port 662 nsew signal input
rlabel metal2 s 101640 99600 101696 100000 6 uP_instr_mem_addr[10]
port 663 nsew signal input
rlabel metal2 s 103488 99600 103544 100000 6 uP_instr_mem_addr[11]
port 664 nsew signal input
rlabel metal2 s 105336 99600 105392 100000 6 uP_instr_mem_addr[12]
port 665 nsew signal input
rlabel metal2 s 81312 99600 81368 100000 6 uP_instr_mem_addr[1]
port 666 nsew signal input
rlabel metal2 s 83776 99600 83832 100000 6 uP_instr_mem_addr[2]
port 667 nsew signal input
rlabel metal2 s 86240 99600 86296 100000 6 uP_instr_mem_addr[3]
port 668 nsew signal input
rlabel metal2 s 88704 99600 88760 100000 6 uP_instr_mem_addr[4]
port 669 nsew signal input
rlabel metal2 s 91168 99600 91224 100000 6 uP_instr_mem_addr[5]
port 670 nsew signal input
rlabel metal2 s 93632 99600 93688 100000 6 uP_instr_mem_addr[6]
port 671 nsew signal input
rlabel metal2 s 96096 99600 96152 100000 6 uP_instr_mem_addr[7]
port 672 nsew signal input
rlabel metal2 s 97944 99600 98000 100000 6 uP_instr_mem_addr[8]
port 673 nsew signal input
rlabel metal2 s 99792 99600 99848 100000 6 uP_instr_mem_addr[9]
port 674 nsew signal input
rlabel metal2 s 79464 99600 79520 100000 6 uP_write_data[0]
port 675 nsew signal input
rlabel metal2 s 102256 99600 102312 100000 6 uP_write_data[10]
port 676 nsew signal input
rlabel metal2 s 104104 99600 104160 100000 6 uP_write_data[11]
port 677 nsew signal input
rlabel metal2 s 105952 99600 106008 100000 6 uP_write_data[12]
port 678 nsew signal input
rlabel metal2 s 107184 99600 107240 100000 6 uP_write_data[13]
port 679 nsew signal input
rlabel metal2 s 108416 99600 108472 100000 6 uP_write_data[14]
port 680 nsew signal input
rlabel metal2 s 109648 99600 109704 100000 6 uP_write_data[15]
port 681 nsew signal input
rlabel metal2 s 81928 99600 81984 100000 6 uP_write_data[1]
port 682 nsew signal input
rlabel metal2 s 84392 99600 84448 100000 6 uP_write_data[2]
port 683 nsew signal input
rlabel metal2 s 86856 99600 86912 100000 6 uP_write_data[3]
port 684 nsew signal input
rlabel metal2 s 89320 99600 89376 100000 6 uP_write_data[4]
port 685 nsew signal input
rlabel metal2 s 91784 99600 91840 100000 6 uP_write_data[5]
port 686 nsew signal input
rlabel metal2 s 94248 99600 94304 100000 6 uP_write_data[6]
port 687 nsew signal input
rlabel metal2 s 96712 99600 96768 100000 6 uP_write_data[7]
port 688 nsew signal input
rlabel metal2 s 98560 99600 98616 100000 6 uP_write_data[8]
port 689 nsew signal input
rlabel metal2 s 100408 99600 100464 100000 6 uP_write_data[9]
port 690 nsew signal input
rlabel metal4 s 2224 1538 2384 98422 6 vdd
port 691 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 98422 6 vdd
port 691 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 98422 6 vdd
port 691 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 98422 6 vdd
port 691 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 98422 6 vdd
port 691 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 98422 6 vdd
port 691 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 98422 6 vdd
port 691 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 98422 6 vdd
port 691 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 98422 6 vdd
port 691 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 98422 6 vdd
port 691 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 98422 6 vdd
port 691 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 98422 6 vdd
port 691 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 98422 6 vss
port 692 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 98422 6 vss
port 692 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 98422 6 vss
port 692 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 98422 6 vss
port 692 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 98422 6 vss
port 692 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 98422 6 vss
port 692 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 98422 6 vss
port 692 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 98422 6 vss
port 692 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 98422 6 vss
port 692 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 98422 6 vss
port 692 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 98422 6 vss
port 692 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 98422 6 vss
port 692 nsew ground bidirectional
rlabel metal2 s 1904 0 1960 400 6 wb_clk_i
port 693 nsew signal input
rlabel metal2 s 2240 0 2296 400 6 wb_rst_i
port 694 nsew signal input
rlabel metal2 s 2576 0 2632 400 6 wbs_ack_o
port 695 nsew signal output
rlabel metal2 s 3920 0 3976 400 6 wbs_adr_i[0]
port 696 nsew signal input
rlabel metal2 s 15344 0 15400 400 6 wbs_adr_i[10]
port 697 nsew signal input
rlabel metal2 s 16352 0 16408 400 6 wbs_adr_i[11]
port 698 nsew signal input
rlabel metal2 s 17360 0 17416 400 6 wbs_adr_i[12]
port 699 nsew signal input
rlabel metal2 s 18368 0 18424 400 6 wbs_adr_i[13]
port 700 nsew signal input
rlabel metal2 s 19376 0 19432 400 6 wbs_adr_i[14]
port 701 nsew signal input
rlabel metal2 s 20384 0 20440 400 6 wbs_adr_i[15]
port 702 nsew signal input
rlabel metal2 s 21392 0 21448 400 6 wbs_adr_i[16]
port 703 nsew signal input
rlabel metal2 s 22400 0 22456 400 6 wbs_adr_i[17]
port 704 nsew signal input
rlabel metal2 s 23408 0 23464 400 6 wbs_adr_i[18]
port 705 nsew signal input
rlabel metal2 s 24416 0 24472 400 6 wbs_adr_i[19]
port 706 nsew signal input
rlabel metal2 s 5264 0 5320 400 6 wbs_adr_i[1]
port 707 nsew signal input
rlabel metal2 s 25424 0 25480 400 6 wbs_adr_i[20]
port 708 nsew signal input
rlabel metal2 s 26432 0 26488 400 6 wbs_adr_i[21]
port 709 nsew signal input
rlabel metal2 s 27440 0 27496 400 6 wbs_adr_i[22]
port 710 nsew signal input
rlabel metal2 s 28448 0 28504 400 6 wbs_adr_i[23]
port 711 nsew signal input
rlabel metal2 s 29456 0 29512 400 6 wbs_adr_i[24]
port 712 nsew signal input
rlabel metal2 s 30464 0 30520 400 6 wbs_adr_i[25]
port 713 nsew signal input
rlabel metal2 s 31472 0 31528 400 6 wbs_adr_i[26]
port 714 nsew signal input
rlabel metal2 s 32480 0 32536 400 6 wbs_adr_i[27]
port 715 nsew signal input
rlabel metal2 s 33488 0 33544 400 6 wbs_adr_i[28]
port 716 nsew signal input
rlabel metal2 s 34496 0 34552 400 6 wbs_adr_i[29]
port 717 nsew signal input
rlabel metal2 s 6608 0 6664 400 6 wbs_adr_i[2]
port 718 nsew signal input
rlabel metal2 s 35504 0 35560 400 6 wbs_adr_i[30]
port 719 nsew signal input
rlabel metal2 s 36512 0 36568 400 6 wbs_adr_i[31]
port 720 nsew signal input
rlabel metal2 s 7952 0 8008 400 6 wbs_adr_i[3]
port 721 nsew signal input
rlabel metal2 s 9296 0 9352 400 6 wbs_adr_i[4]
port 722 nsew signal input
rlabel metal2 s 10304 0 10360 400 6 wbs_adr_i[5]
port 723 nsew signal input
rlabel metal2 s 11312 0 11368 400 6 wbs_adr_i[6]
port 724 nsew signal input
rlabel metal2 s 12320 0 12376 400 6 wbs_adr_i[7]
port 725 nsew signal input
rlabel metal2 s 13328 0 13384 400 6 wbs_adr_i[8]
port 726 nsew signal input
rlabel metal2 s 14336 0 14392 400 6 wbs_adr_i[9]
port 727 nsew signal input
rlabel metal2 s 2912 0 2968 400 6 wbs_cyc_i
port 728 nsew signal input
rlabel metal2 s 4256 0 4312 400 6 wbs_dat_i[0]
port 729 nsew signal input
rlabel metal2 s 15680 0 15736 400 6 wbs_dat_i[10]
port 730 nsew signal input
rlabel metal2 s 16688 0 16744 400 6 wbs_dat_i[11]
port 731 nsew signal input
rlabel metal2 s 17696 0 17752 400 6 wbs_dat_i[12]
port 732 nsew signal input
rlabel metal2 s 18704 0 18760 400 6 wbs_dat_i[13]
port 733 nsew signal input
rlabel metal2 s 19712 0 19768 400 6 wbs_dat_i[14]
port 734 nsew signal input
rlabel metal2 s 20720 0 20776 400 6 wbs_dat_i[15]
port 735 nsew signal input
rlabel metal2 s 21728 0 21784 400 6 wbs_dat_i[16]
port 736 nsew signal input
rlabel metal2 s 22736 0 22792 400 6 wbs_dat_i[17]
port 737 nsew signal input
rlabel metal2 s 23744 0 23800 400 6 wbs_dat_i[18]
port 738 nsew signal input
rlabel metal2 s 24752 0 24808 400 6 wbs_dat_i[19]
port 739 nsew signal input
rlabel metal2 s 5600 0 5656 400 6 wbs_dat_i[1]
port 740 nsew signal input
rlabel metal2 s 25760 0 25816 400 6 wbs_dat_i[20]
port 741 nsew signal input
rlabel metal2 s 26768 0 26824 400 6 wbs_dat_i[21]
port 742 nsew signal input
rlabel metal2 s 27776 0 27832 400 6 wbs_dat_i[22]
port 743 nsew signal input
rlabel metal2 s 28784 0 28840 400 6 wbs_dat_i[23]
port 744 nsew signal input
rlabel metal2 s 29792 0 29848 400 6 wbs_dat_i[24]
port 745 nsew signal input
rlabel metal2 s 30800 0 30856 400 6 wbs_dat_i[25]
port 746 nsew signal input
rlabel metal2 s 31808 0 31864 400 6 wbs_dat_i[26]
port 747 nsew signal input
rlabel metal2 s 32816 0 32872 400 6 wbs_dat_i[27]
port 748 nsew signal input
rlabel metal2 s 33824 0 33880 400 6 wbs_dat_i[28]
port 749 nsew signal input
rlabel metal2 s 34832 0 34888 400 6 wbs_dat_i[29]
port 750 nsew signal input
rlabel metal2 s 6944 0 7000 400 6 wbs_dat_i[2]
port 751 nsew signal input
rlabel metal2 s 35840 0 35896 400 6 wbs_dat_i[30]
port 752 nsew signal input
rlabel metal2 s 36848 0 36904 400 6 wbs_dat_i[31]
port 753 nsew signal input
rlabel metal2 s 8288 0 8344 400 6 wbs_dat_i[3]
port 754 nsew signal input
rlabel metal2 s 9632 0 9688 400 6 wbs_dat_i[4]
port 755 nsew signal input
rlabel metal2 s 10640 0 10696 400 6 wbs_dat_i[5]
port 756 nsew signal input
rlabel metal2 s 11648 0 11704 400 6 wbs_dat_i[6]
port 757 nsew signal input
rlabel metal2 s 12656 0 12712 400 6 wbs_dat_i[7]
port 758 nsew signal input
rlabel metal2 s 13664 0 13720 400 6 wbs_dat_i[8]
port 759 nsew signal input
rlabel metal2 s 14672 0 14728 400 6 wbs_dat_i[9]
port 760 nsew signal input
rlabel metal2 s 4592 0 4648 400 6 wbs_dat_o[0]
port 761 nsew signal output
rlabel metal2 s 16016 0 16072 400 6 wbs_dat_o[10]
port 762 nsew signal output
rlabel metal2 s 17024 0 17080 400 6 wbs_dat_o[11]
port 763 nsew signal output
rlabel metal2 s 18032 0 18088 400 6 wbs_dat_o[12]
port 764 nsew signal output
rlabel metal2 s 19040 0 19096 400 6 wbs_dat_o[13]
port 765 nsew signal output
rlabel metal2 s 20048 0 20104 400 6 wbs_dat_o[14]
port 766 nsew signal output
rlabel metal2 s 21056 0 21112 400 6 wbs_dat_o[15]
port 767 nsew signal output
rlabel metal2 s 22064 0 22120 400 6 wbs_dat_o[16]
port 768 nsew signal output
rlabel metal2 s 23072 0 23128 400 6 wbs_dat_o[17]
port 769 nsew signal output
rlabel metal2 s 24080 0 24136 400 6 wbs_dat_o[18]
port 770 nsew signal output
rlabel metal2 s 25088 0 25144 400 6 wbs_dat_o[19]
port 771 nsew signal output
rlabel metal2 s 5936 0 5992 400 6 wbs_dat_o[1]
port 772 nsew signal output
rlabel metal2 s 26096 0 26152 400 6 wbs_dat_o[20]
port 773 nsew signal output
rlabel metal2 s 27104 0 27160 400 6 wbs_dat_o[21]
port 774 nsew signal output
rlabel metal2 s 28112 0 28168 400 6 wbs_dat_o[22]
port 775 nsew signal output
rlabel metal2 s 29120 0 29176 400 6 wbs_dat_o[23]
port 776 nsew signal output
rlabel metal2 s 30128 0 30184 400 6 wbs_dat_o[24]
port 777 nsew signal output
rlabel metal2 s 31136 0 31192 400 6 wbs_dat_o[25]
port 778 nsew signal output
rlabel metal2 s 32144 0 32200 400 6 wbs_dat_o[26]
port 779 nsew signal output
rlabel metal2 s 33152 0 33208 400 6 wbs_dat_o[27]
port 780 nsew signal output
rlabel metal2 s 34160 0 34216 400 6 wbs_dat_o[28]
port 781 nsew signal output
rlabel metal2 s 35168 0 35224 400 6 wbs_dat_o[29]
port 782 nsew signal output
rlabel metal2 s 7280 0 7336 400 6 wbs_dat_o[2]
port 783 nsew signal output
rlabel metal2 s 36176 0 36232 400 6 wbs_dat_o[30]
port 784 nsew signal output
rlabel metal2 s 37184 0 37240 400 6 wbs_dat_o[31]
port 785 nsew signal output
rlabel metal2 s 8624 0 8680 400 6 wbs_dat_o[3]
port 786 nsew signal output
rlabel metal2 s 9968 0 10024 400 6 wbs_dat_o[4]
port 787 nsew signal output
rlabel metal2 s 10976 0 11032 400 6 wbs_dat_o[5]
port 788 nsew signal output
rlabel metal2 s 11984 0 12040 400 6 wbs_dat_o[6]
port 789 nsew signal output
rlabel metal2 s 12992 0 13048 400 6 wbs_dat_o[7]
port 790 nsew signal output
rlabel metal2 s 14000 0 14056 400 6 wbs_dat_o[8]
port 791 nsew signal output
rlabel metal2 s 15008 0 15064 400 6 wbs_dat_o[9]
port 792 nsew signal output
rlabel metal2 s 4928 0 4984 400 6 wbs_sel_i[0]
port 793 nsew signal input
rlabel metal2 s 6272 0 6328 400 6 wbs_sel_i[1]
port 794 nsew signal input
rlabel metal2 s 7616 0 7672 400 6 wbs_sel_i[2]
port 795 nsew signal input
rlabel metal2 s 8960 0 9016 400 6 wbs_sel_i[3]
port 796 nsew signal input
rlabel metal2 s 3248 0 3304 400 6 wbs_stb_i
port 797 nsew signal input
rlabel metal2 s 3584 0 3640 400 6 wbs_we_i
port 798 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 180000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8730786
string GDS_FILE /home/radhe/tapeout_projects/gf_new/sathvik/openlane/io_interface/runs/22_12_10_14_28/results/signoff/io_interface.magic.gds
string GDS_START 171848
<< end >>

