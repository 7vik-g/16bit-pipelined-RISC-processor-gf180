// This is the unpowered netlist.
module processor (Dataw_en,
    Serial_input,
    Serial_output,
    clk,
    hlt,
    reset,
    start,
    data_mem_addr,
    instr,
    instr_mem_addr,
    read_data,
    write_data);
 output Dataw_en;
 input Serial_input;
 output Serial_output;
 input clk;
 output hlt;
 input reset;
 input start;
 output [7:0] data_mem_addr;
 input [15:0] instr;
 output [12:0] instr_mem_addr;
 input [15:0] read_data;
 output [15:0] write_data;

 wire \Arithmetic_Logic_Unit.ALU_000.ALU_func[0] ;
 wire \Arithmetic_Logic_Unit.ALU_000.ALU_func[1] ;
 wire \Arithmetic_Logic_Unit.ALU_000.ALU_func[2] ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[0].i2 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[0].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i0 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i2 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[11].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[12].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[13].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[14].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[1].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[2].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[3].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[4].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[6].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.Y_CY[7].i3 ;
 wire \Arithmetic_Logic_Unit.ALU_001.p_Z ;
 wire \Arithmetic_Logic_Unit.op ;
 wire \Control_unit1.instr_decoder1.A[0] ;
 wire \Control_unit1.instr_decoder1.A[1] ;
 wire \Control_unit1.instr_decoder1.A[2] ;
 wire \Control_unit1.instr_stage1[0] ;
 wire \Control_unit1.instr_stage1[10] ;
 wire \Control_unit1.instr_stage1[11] ;
 wire \Control_unit1.instr_stage1[12] ;
 wire \Control_unit1.instr_stage1[1] ;
 wire \Control_unit1.instr_stage1[2] ;
 wire \Control_unit1.instr_stage1[3] ;
 wire \Control_unit1.instr_stage1[4] ;
 wire \Control_unit1.instr_stage1[5] ;
 wire \Control_unit1.instr_stage1[6] ;
 wire \Control_unit1.instr_stage1[7] ;
 wire \Control_unit1.instr_stage1[8] ;
 wire \Control_unit1.instr_stage1[9] ;
 wire \Control_unit2.instr_decoder2.A[1] ;
 wire \Control_unit2.instr_decoder2.A[2] ;
 wire \Control_unit2.instr_stage2[10] ;
 wire \Control_unit2.instr_stage2[11] ;
 wire \Control_unit2.instr_stage2[12] ;
 wire \Control_unit2.instr_stage2[3] ;
 wire \Control_unit2.instr_stage2[4] ;
 wire \Control_unit2.instr_stage2[5] ;
 wire \Control_unit2.instr_stage2[6] ;
 wire \Control_unit2.instr_stage2[7] ;
 wire \Control_unit2.instr_stage2[8] ;
 wire \Control_unit2.instr_stage2[9] ;
 wire \Stack_pointer.SP[0] ;
 wire \Stack_pointer.SP[1] ;
 wire \Stack_pointer.SP[2] ;
 wire \Stack_pointer.SP[3] ;
 wire \Stack_pointer.SP[4] ;
 wire \Stack_pointer.SP[5] ;
 wire \Stack_pointer.SP[6] ;
 wire \Stack_pointer.SP[7] ;
 wire \Stack_pointer.SP_next[0] ;
 wire \Stack_pointer.SP_next[1] ;
 wire \Stack_pointer.SP_next[2] ;
 wire \Stack_pointer.SP_next[3] ;
 wire \Stack_pointer.SP_next[4] ;
 wire \Stack_pointer.SP_next[5] ;
 wire \Stack_pointer.SP_next[6] ;
 wire \Stack_pointer.SP_next[7] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;

 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2382_ (.I(\Arithmetic_Logic_Unit.ALU_000.ALU_func[0] ),
    .Z(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2383_ (.I(_2078_),
    .Z(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2384_ (.I(\Arithmetic_Logic_Unit.ALU_000.ALU_func[2] ),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2385_ (.I(\Arithmetic_Logic_Unit.ALU_000.ALU_func[1] ),
    .Z(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2386_ (.I(_2081_),
    .Z(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2387_ (.I(_2082_),
    .Z(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2388_ (.I(_2083_),
    .Z(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2389_ (.I(\Control_unit2.instr_decoder2.A[2] ),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2390_ (.A1(\Arithmetic_Logic_Unit.op ),
    .A2(_2085_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2391_ (.A1(_2080_),
    .A2(\Control_unit2.instr_decoder2.A[1] ),
    .A3(_2084_),
    .A4(_2086_),
    .ZN(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2392_ (.A1(_2079_),
    .A2(_2087_),
    .ZN(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2393_ (.I(\Control_unit2.instr_stage2[12] ),
    .Z(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2394_ (.A1(_2089_),
    .A2(\Control_unit2.instr_stage2[11] ),
    .ZN(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2395_ (.A1(_2088_),
    .A2(_2090_),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2396_ (.I(_2091_),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2397_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[0].i3 ),
    .Z(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2398_ (.A1(\Arithmetic_Logic_Unit.ALU_000.ALU_func[0] ),
    .A2(\Arithmetic_Logic_Unit.ALU_000.ALU_func[1] ),
    .Z(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2399_ (.A1(_2080_),
    .A2(_2093_),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2400_ (.I(_2094_),
    .Z(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2401_ (.I(_2095_),
    .Z(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2402_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[0].i3 ),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2403_ (.A1(_2078_),
    .A2(_2081_),
    .B(\Arithmetic_Logic_Unit.ALU_000.ALU_func[2] ),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2404_ (.I(_2098_),
    .Z(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2405_ (.A1(_2083_),
    .A2(_2097_),
    .B(_2099_),
    .ZN(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2406_ (.I(\Arithmetic_Logic_Unit.ALU_000.ALU_func[2] ),
    .Z(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2407_ (.I(_2081_),
    .ZN(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2408_ (.A1(_2101_),
    .A2(_2102_),
    .B(_2093_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2409_ (.I(_2103_),
    .Z(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2410_ (.A1(_2092_),
    .A2(_2096_),
    .A3(_2100_),
    .A4(_2104_),
    .Z(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2411_ (.I(_2092_),
    .Z(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2412_ (.I(_2094_),
    .Z(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2413_ (.I(_2107_),
    .Z(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2414_ (.I0(\Arithmetic_Logic_Unit.ALU_000.ALU_func[2] ),
    .I1(_2078_),
    .S(_2081_),
    .Z(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2415_ (.I(_2109_),
    .Z(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2416_ (.A1(_2092_),
    .A2(_2110_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2417_ (.A1(_2106_),
    .A2(_2108_),
    .B1(_2100_),
    .B2(_2111_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2418_ (.A1(_2105_),
    .A2(_2112_),
    .Z(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2419_ (.I(\Control_unit1.instr_decoder1.A[0] ),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2420_ (.A1(\Control_unit1.instr_decoder1.A[2] ),
    .A2(\Control_unit1.instr_decoder1.A[1] ),
    .Z(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2421_ (.A1(\Control_unit1.instr_stage1[3] ),
    .A2(\Control_unit1.instr_stage1[1] ),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2422_ (.A1(_2114_),
    .A2(\Control_unit1.instr_stage1[2] ),
    .A3(_2115_),
    .A4(_2116_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2423_ (.I0(net37),
    .I1(net1),
    .S(_2117_),
    .Z(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _2424_ (.I(_2079_),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2425_ (.A1(_2083_),
    .A2(_2118_),
    .B(_2119_),
    .C(_2101_),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2426_ (.I(net37),
    .ZN(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2427_ (.I(net1),
    .ZN(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2428_ (.I0(_2121_),
    .I1(_2122_),
    .S(_2117_),
    .Z(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2429_ (.I(_2102_),
    .Z(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2430_ (.A1(_2078_),
    .A2(_2124_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2431_ (.I(_2125_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2432_ (.A1(_2079_),
    .A2(_2123_),
    .B(_2126_),
    .C(_2080_),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2433_ (.A1(_2120_),
    .A2(_2127_),
    .Z(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2434_ (.A1(_2113_),
    .A2(_2128_),
    .Z(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2435_ (.I(_2102_),
    .Z(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2436_ (.I(_2130_),
    .Z(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2437_ (.I(_2131_),
    .Z(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2438_ (.I(_2132_),
    .Z(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2439_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[1].i3 ),
    .Z(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2440_ (.I(_2134_),
    .Z(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2441_ (.I(_2093_),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2442_ (.I(_2136_),
    .Z(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2443_ (.I(_2125_),
    .Z(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2444_ (.I(_2138_),
    .Z(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2445_ (.A1(_2133_),
    .A2(_2106_),
    .B1(_2135_),
    .B2(_2137_),
    .C1(_2139_),
    .C2(_2118_),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2446_ (.I(\Arithmetic_Logic_Unit.op ),
    .Z(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2447_ (.I(_2141_),
    .Z(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2448_ (.I(_2142_),
    .Z(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2449_ (.I0(_2129_),
    .I1(_2140_),
    .S(_2143_),
    .Z(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2450_ (.I(_2144_),
    .Z(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2451_ (.I(_2145_),
    .Z(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2452_ (.I(_2146_),
    .ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2453_ (.I(_2141_),
    .Z(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2454_ (.I(_2147_),
    .Z(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2455_ (.I(_2095_),
    .Z(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2456_ (.I(_2103_),
    .Z(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2457_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[1].i3 ),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2458_ (.I(_2098_),
    .Z(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2459_ (.A1(_2082_),
    .A2(_2151_),
    .B(_2152_),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _2460_ (.A1(_2134_),
    .A2(_2149_),
    .A3(_2150_),
    .A4(_2153_),
    .Z(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2461_ (.I(_2109_),
    .Z(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2462_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[1].i3 ),
    .A2(_2155_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2463_ (.A1(_2134_),
    .A2(_2096_),
    .B1(_2156_),
    .B2(_2153_),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2464_ (.A1(_2154_),
    .A2(_2157_),
    .Z(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2465_ (.I(_2112_),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2466_ (.A1(_2159_),
    .A2(_2128_),
    .B(_2105_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2467_ (.A1(_2158_),
    .A2(_2160_),
    .Z(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2468_ (.I(_2142_),
    .Z(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2469_ (.I(_2132_),
    .Z(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2470_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[2].i3 ),
    .Z(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2471_ (.I(_2164_),
    .Z(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2472_ (.I(_2136_),
    .Z(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2473_ (.I(_2166_),
    .Z(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2474_ (.A1(_2163_),
    .A2(_2135_),
    .B1(_2165_),
    .B2(_2167_),
    .C1(_2139_),
    .C2(_2106_),
    .ZN(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2475_ (.A1(_2162_),
    .A2(_2168_),
    .ZN(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2476_ (.A1(_2148_),
    .A2(_2161_),
    .B(_2169_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2477_ (.I(_2170_),
    .Z(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2478_ (.I(_2171_),
    .Z(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2479_ (.I(_2172_),
    .ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2480_ (.A1(_2113_),
    .A2(_2158_),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2481_ (.A1(_2092_),
    .A2(_2096_),
    .A3(_2100_),
    .A4(_2104_),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2482_ (.A1(_2174_),
    .A2(_2154_),
    .A3(_2157_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2483_ (.A1(_2128_),
    .A2(_2173_),
    .B(_2175_),
    .C(_2154_),
    .ZN(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2484_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[2].i3 ),
    .ZN(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2485_ (.A1(_2082_),
    .A2(_2177_),
    .B(_2099_),
    .ZN(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2486_ (.A1(_2164_),
    .A2(_2149_),
    .A3(_2150_),
    .A4(_2178_),
    .Z(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2487_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[2].i3 ),
    .A2(_2110_),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2488_ (.A1(_2164_),
    .A2(_2096_),
    .B1(_2180_),
    .B2(_2178_),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2489_ (.A1(_2179_),
    .A2(_2181_),
    .Z(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2490_ (.A1(_2176_),
    .A2(_2182_),
    .Z(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2491_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[3].i3 ),
    .Z(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2492_ (.I(_2184_),
    .Z(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2493_ (.A1(_2163_),
    .A2(_2165_),
    .B1(_2185_),
    .B2(_2167_),
    .C1(_2139_),
    .C2(_2135_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2494_ (.A1(_2162_),
    .A2(_2186_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2495_ (.A1(_2148_),
    .A2(_2183_),
    .B(_2187_),
    .ZN(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2496_ (.I(_2188_),
    .Z(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2497_ (.I(_2189_),
    .Z(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2498_ (.I(_2190_),
    .ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2499_ (.I(_2107_),
    .Z(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2500_ (.A1(_2184_),
    .A2(_2110_),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2501_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[3].i3 ),
    .ZN(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2502_ (.A1(_2082_),
    .A2(_2193_),
    .B(_2098_),
    .ZN(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _2503_ (.A1(_2184_),
    .A2(_2191_),
    .B1(_2192_),
    .B2(_2194_),
    .ZN(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2504_ (.A1(_2184_),
    .A2(_2107_),
    .A3(_2150_),
    .A4(_2194_),
    .Z(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2505_ (.I(_2196_),
    .Z(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2506_ (.A1(_2195_),
    .A2(_2197_),
    .ZN(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2507_ (.A1(_2128_),
    .A2(_2173_),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2508_ (.A1(_2134_),
    .A2(_2191_),
    .A3(_2104_),
    .A4(_2153_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2509_ (.A1(_2200_),
    .A2(_2179_),
    .A3(_2181_),
    .ZN(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2510_ (.A1(_2175_),
    .A2(_2179_),
    .A3(_2201_),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2511_ (.A1(_2199_),
    .A2(_2182_),
    .B(_2202_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2512_ (.A1(_2198_),
    .A2(_2203_),
    .ZN(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2513_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[4].i3 ),
    .Z(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2514_ (.I(_2205_),
    .Z(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2515_ (.I(_2166_),
    .Z(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2516_ (.I(_2138_),
    .Z(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2517_ (.A1(_2163_),
    .A2(_2185_),
    .B1(_2206_),
    .B2(_2207_),
    .C1(_2208_),
    .C2(_2165_),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2518_ (.I0(_2204_),
    .I1(_2209_),
    .S(_2162_),
    .Z(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2519_ (.I(_2210_),
    .Z(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2520_ (.I(_2211_),
    .Z(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2521_ (.I(_2212_),
    .ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2522_ (.A1(_2154_),
    .A2(_2157_),
    .A3(_2179_),
    .A4(_2181_),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2523_ (.A1(_2105_),
    .A2(_2112_),
    .A3(_2195_),
    .A4(_2197_),
    .ZN(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2524_ (.A1(_2120_),
    .A2(_2127_),
    .A3(_2213_),
    .A4(_2214_),
    .Z(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2525_ (.A1(_2164_),
    .A2(_2108_),
    .A3(_2104_),
    .A4(_2178_),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2526_ (.A1(_2216_),
    .A2(_2195_),
    .A3(_2196_),
    .ZN(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2527_ (.A1(_2175_),
    .A2(_2197_),
    .A3(_2201_),
    .A4(_2217_),
    .Z(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2528_ (.A1(_2205_),
    .A2(_2149_),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2529_ (.A1(_2130_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[4].i3 ),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2530_ (.A1(_2205_),
    .A2(_2155_),
    .B1(_2220_),
    .B2(_2099_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2531_ (.A1(_2219_),
    .A2(_2221_),
    .Z(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2532_ (.I(_2222_),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2533_ (.A1(_2215_),
    .A2(_2218_),
    .B(_2223_),
    .ZN(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _2534_ (.A1(_2120_),
    .A2(_2127_),
    .A3(_2213_),
    .A4(_2214_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2535_ (.A1(_2175_),
    .A2(_2197_),
    .A3(_2201_),
    .A4(_2217_),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2536_ (.A1(_2225_),
    .A2(_2226_),
    .A3(_2222_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2537_ (.A1(_2224_),
    .A2(_2227_),
    .Z(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2538_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ),
    .Z(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2539_ (.A1(_2229_),
    .A2(_2166_),
    .B1(_2138_),
    .B2(_2185_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2540_ (.A1(_2142_),
    .A2(_2220_),
    .A3(_2230_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2541_ (.A1(_2147_),
    .A2(_2228_),
    .B(_2231_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2542_ (.I(_2232_),
    .ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2543_ (.I(_2162_),
    .Z(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2544_ (.I(_2107_),
    .Z(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2545_ (.A1(_2205_),
    .A2(_2234_),
    .A3(_2221_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2546_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ),
    .A2(_2095_),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2547_ (.A1(_2130_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2548_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ),
    .A2(_2109_),
    .B1(_2237_),
    .B2(_2152_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2549_ (.A1(_2236_),
    .A2(_2238_),
    .Z(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2550_ (.I(_2239_),
    .Z(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2551_ (.A1(_2235_),
    .A2(_2224_),
    .A3(_2240_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2552_ (.A1(_2222_),
    .A2(_2239_),
    .Z(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2553_ (.A1(_2225_),
    .A2(_2226_),
    .B(_2242_),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2554_ (.A1(_2235_),
    .A2(_2240_),
    .ZN(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2555_ (.I(_2244_),
    .Z(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2556_ (.A1(_2243_),
    .A2(_2245_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2557_ (.A1(_2241_),
    .A2(_2246_),
    .Z(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2558_ (.I(_2143_),
    .Z(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2559_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[6].i3 ),
    .Z(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2560_ (.I(_2249_),
    .Z(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2561_ (.I(_2137_),
    .Z(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2562_ (.I(_2125_),
    .Z(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2563_ (.I(_2252_),
    .Z(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2564_ (.A1(_2250_),
    .A2(_2251_),
    .B1(_2253_),
    .B2(_2206_),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2565_ (.A1(_2248_),
    .A2(_2237_),
    .A3(_2254_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2566_ (.A1(_2233_),
    .A2(_2247_),
    .B(_2255_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2567_ (.I(_2256_),
    .Z(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2568_ (.I(_2257_),
    .ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2569_ (.I(_2143_),
    .Z(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2570_ (.I(_2108_),
    .Z(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2571_ (.I(_2259_),
    .Z(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2572_ (.I(_2260_),
    .Z(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2573_ (.A1(_2229_),
    .A2(_2261_),
    .A3(_2238_),
    .Z(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2574_ (.A1(_2249_),
    .A2(_2095_),
    .ZN(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2575_ (.A1(_2130_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[6].i3 ),
    .ZN(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2576_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[6].i3 ),
    .A2(_2155_),
    .B1(_2264_),
    .B2(_2152_),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2577_ (.A1(_2263_),
    .A2(_2265_),
    .Z(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2578_ (.I(_2266_),
    .Z(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2579_ (.I(_2267_),
    .ZN(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2580_ (.A1(_2262_),
    .A2(_2243_),
    .A3(_2245_),
    .A4(_2268_),
    .Z(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2581_ (.A1(_2262_),
    .A2(_2243_),
    .A3(_2245_),
    .B(_2268_),
    .ZN(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2582_ (.A1(_2269_),
    .A2(_2270_),
    .Z(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2583_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[7].i3 ),
    .Z(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2584_ (.I(_2272_),
    .Z(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2585_ (.I(_2229_),
    .Z(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2586_ (.A1(_2273_),
    .A2(_2251_),
    .B1(_2253_),
    .B2(_2274_),
    .ZN(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2587_ (.A1(_2148_),
    .A2(_2264_),
    .A3(_2275_),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2588_ (.A1(_2258_),
    .A2(_2271_),
    .B(_2276_),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2589_ (.I(_2277_),
    .Z(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2590_ (.I(_2278_),
    .ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2591_ (.I(_2147_),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2592_ (.I(_2279_),
    .Z(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2593_ (.A1(_2124_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[7].i3 ),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2594_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i2 ),
    .Z(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2595_ (.I(_2282_),
    .Z(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2596_ (.A1(_2283_),
    .A2(_2167_),
    .B1(_2139_),
    .B2(_2249_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2597_ (.A1(_2281_),
    .A2(_2284_),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2598_ (.A1(_2272_),
    .A2(_2149_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2599_ (.A1(_2272_),
    .A2(_2110_),
    .B1(_2281_),
    .B2(_2099_),
    .ZN(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2600_ (.A1(_2286_),
    .A2(_2287_),
    .Z(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2601_ (.A1(_2249_),
    .A2(_2259_),
    .A3(_2265_),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2602_ (.I(_2289_),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2603_ (.A1(_2229_),
    .A2(_2234_),
    .A3(_2238_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2604_ (.A1(_2291_),
    .A2(_2267_),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2605_ (.A1(_2245_),
    .A2(_2290_),
    .A3(_2292_),
    .ZN(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2606_ (.A1(_2224_),
    .A2(_2240_),
    .A3(_2267_),
    .B(_2293_),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2607_ (.A1(_2288_),
    .A2(_2294_),
    .Z(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2608_ (.A1(_2280_),
    .A2(_2295_),
    .ZN(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2609_ (.A1(_2280_),
    .A2(_2285_),
    .B(_2296_),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2610_ (.I(_2297_),
    .Z(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2611_ (.I(_2298_),
    .ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2612_ (.A1(_2222_),
    .A2(_2240_),
    .A3(_2267_),
    .A4(_2288_),
    .ZN(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2613_ (.A1(_2215_),
    .A2(_2218_),
    .B(_2299_),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2614_ (.A1(_2272_),
    .A2(_2259_),
    .A3(_2287_),
    .Z(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2615_ (.A1(_2289_),
    .A2(_2288_),
    .ZN(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2616_ (.A1(_2244_),
    .A2(_2301_),
    .A3(_2292_),
    .A4(_2302_),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2617_ (.A1(_2282_),
    .A2(_2234_),
    .ZN(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2618_ (.I(_2155_),
    .Z(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2619_ (.A1(_2131_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i2 ),
    .ZN(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2620_ (.I(_2152_),
    .Z(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2621_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i2 ),
    .A2(_2305_),
    .B1(_2306_),
    .B2(_2307_),
    .ZN(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2622_ (.A1(_2304_),
    .A2(_2308_),
    .Z(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2623_ (.A1(_2300_),
    .A2(_2303_),
    .B(_2309_),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2624_ (.A1(_2266_),
    .A2(_2288_),
    .Z(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2625_ (.A1(_2225_),
    .A2(_2226_),
    .B(_2242_),
    .C(_2311_),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _2626_ (.A1(_2244_),
    .A2(_2301_),
    .A3(_2292_),
    .A4(_2302_),
    .Z(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2627_ (.A1(_2304_),
    .A2(_2308_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2628_ (.A1(_2312_),
    .A2(_2313_),
    .A3(_2314_),
    .ZN(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2629_ (.A1(_2310_),
    .A2(_2315_),
    .B(_2280_),
    .ZN(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2630_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i0 ),
    .Z(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2631_ (.I(_2317_),
    .Z(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2632_ (.A1(_2133_),
    .A2(_2283_),
    .B1(_2318_),
    .B2(_2137_),
    .C1(_2252_),
    .C2(_2273_),
    .ZN(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2633_ (.A1(_2258_),
    .A2(_2319_),
    .ZN(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2634_ (.A1(_2316_),
    .A2(_2320_),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2635_ (.I(_2321_),
    .Z(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2636_ (.I(_2322_),
    .ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2637_ (.A1(_2282_),
    .A2(_2259_),
    .A3(_2308_),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2638_ (.A1(_2317_),
    .A2(_2191_),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2639_ (.A1(_2124_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i0 ),
    .ZN(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2640_ (.A1(_2317_),
    .A2(_2305_),
    .B1(_2325_),
    .B2(_2307_),
    .ZN(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2641_ (.A1(_2324_),
    .A2(_2326_),
    .Z(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2642_ (.A1(_2323_),
    .A2(_2327_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2643_ (.A1(_2309_),
    .A2(_2327_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2644_ (.A1(_2312_),
    .A2(_2313_),
    .B(_2329_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2645_ (.A1(_2323_),
    .A2(_2327_),
    .Z(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2646_ (.A1(_2310_),
    .A2(_2328_),
    .B(_2330_),
    .C(_2331_),
    .ZN(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2647_ (.A1(_2133_),
    .A2(_2318_),
    .B1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ),
    .B2(_2166_),
    .C1(_2252_),
    .C2(_2282_),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2648_ (.I0(_2332_),
    .I1(_2333_),
    .S(_2143_),
    .Z(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2649_ (.I(_2334_),
    .Z(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2650_ (.I(_2335_),
    .Z(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2651_ (.I(_2336_),
    .ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2652_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[11].i3 ),
    .Z(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2653_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ),
    .ZN(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2654_ (.A1(_2083_),
    .A2(_2338_),
    .ZN(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2655_ (.A1(_2337_),
    .A2(_2137_),
    .B1(_2252_),
    .B2(_2318_),
    .C(_2339_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2656_ (.A1(_2248_),
    .A2(_2340_),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2657_ (.I(_2234_),
    .Z(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2658_ (.A1(_2317_),
    .A2(_2342_),
    .A3(_2326_),
    .ZN(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2659_ (.A1(_2343_),
    .A2(_2331_),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2660_ (.I(_2344_),
    .ZN(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2661_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ),
    .A2(_2191_),
    .ZN(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2662_ (.A1(_2101_),
    .A2(_2136_),
    .A3(_2339_),
    .B1(_2150_),
    .B2(_2338_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2663_ (.A1(_2346_),
    .A2(_2347_),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2664_ (.A1(_2330_),
    .A2(_2345_),
    .B(_2348_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2665_ (.A1(_2300_),
    .A2(_2303_),
    .B(_2309_),
    .C(_2327_),
    .ZN(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2666_ (.I(_2348_),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2667_ (.A1(_2350_),
    .A2(_2351_),
    .A3(_2344_),
    .ZN(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2668_ (.A1(_2349_),
    .A2(_2352_),
    .B(_2280_),
    .ZN(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2669_ (.A1(_2341_),
    .A2(_2353_),
    .ZN(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2670_ (.I(_2354_),
    .Z(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2671_ (.I(_2355_),
    .ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2672_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[11].i3 ),
    .A2(_2108_),
    .ZN(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2673_ (.A1(_2124_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[11].i3 ),
    .ZN(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2674_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[11].i3 ),
    .A2(_2305_),
    .B1(_2357_),
    .B2(_2307_),
    .ZN(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2675_ (.A1(_2356_),
    .A2(_2358_),
    .Z(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2676_ (.A1(_2346_),
    .A2(_2347_),
    .Z(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2677_ (.A1(_2343_),
    .A2(_2348_),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2678_ (.A1(_2331_),
    .A2(_2360_),
    .A3(_2361_),
    .ZN(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2679_ (.A1(_2350_),
    .A2(_2351_),
    .B(_2362_),
    .ZN(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2680_ (.A1(_2359_),
    .A2(_2363_),
    .Z(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2681_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[12].i3 ),
    .Z(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2682_ (.I(_2365_),
    .Z(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2683_ (.I(_2357_),
    .ZN(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2684_ (.A1(_2366_),
    .A2(_2136_),
    .B1(_2138_),
    .B2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ),
    .C(_2367_),
    .ZN(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2685_ (.A1(_2142_),
    .A2(_2368_),
    .ZN(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2686_ (.A1(_2147_),
    .A2(_2364_),
    .B(_2369_),
    .ZN(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2687_ (.I(_2370_),
    .ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2688_ (.A1(_2365_),
    .A2(_2342_),
    .ZN(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2689_ (.I(_2305_),
    .Z(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2690_ (.A1(_2131_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[12].i3 ),
    .ZN(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2691_ (.I(_2307_),
    .Z(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2692_ (.A1(_2365_),
    .A2(_2372_),
    .B1(_2373_),
    .B2(_2374_),
    .ZN(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2693_ (.A1(_2371_),
    .A2(_2375_),
    .Z(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2694_ (.I(_2376_),
    .ZN(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2695_ (.A1(_2348_),
    .A2(_2359_),
    .ZN(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2696_ (.A1(_2329_),
    .A2(_2378_),
    .ZN(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2697_ (.A1(_2300_),
    .A2(_2303_),
    .B(_2379_),
    .ZN(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2698_ (.A1(_2337_),
    .A2(_2260_),
    .A3(_2358_),
    .ZN(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2699_ (.A1(_2360_),
    .A2(_2359_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2700_ (.A1(_2331_),
    .A2(_2381_),
    .A3(_2361_),
    .A4(_0559_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2701_ (.A1(_2377_),
    .A2(_2380_),
    .A3(_0560_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2702_ (.A1(_2312_),
    .A2(_2313_),
    .B(_2329_),
    .C(_2378_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2703_ (.I(_0560_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2704_ (.A1(_0562_),
    .A2(_0563_),
    .B(_2376_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2705_ (.A1(_0561_),
    .A2(_0564_),
    .B(_2279_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2706_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[13].i3 ),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2707_ (.I(_0566_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2708_ (.A1(_2163_),
    .A2(_2366_),
    .B1(_0567_),
    .B2(_2167_),
    .C1(_2208_),
    .C2(_2337_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2709_ (.A1(_2148_),
    .A2(_0568_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2710_ (.A1(_0565_),
    .A2(_0569_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2711_ (.I(_0570_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2712_ (.I(_0571_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2713_ (.I(_0572_),
    .ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2714_ (.A1(_2380_),
    .A2(_0560_),
    .B(_2377_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2715_ (.A1(_2365_),
    .A2(_2261_),
    .A3(_2375_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2716_ (.A1(_2131_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[13].i3 ),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2717_ (.A1(_0566_),
    .A2(_2372_),
    .B1(_0575_),
    .B2(_2374_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2718_ (.A1(_0566_),
    .A2(_2342_),
    .A3(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2719_ (.I(_0577_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2720_ (.A1(_0566_),
    .A2(_2342_),
    .B(_0576_),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2721_ (.A1(_0578_),
    .A2(_0579_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2722_ (.A1(_0574_),
    .A2(_0580_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2723_ (.A1(_2376_),
    .A2(_0580_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2724_ (.A1(_0562_),
    .A2(_0563_),
    .B(_0582_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2725_ (.A1(_0574_),
    .A2(_0580_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2726_ (.A1(_0573_),
    .A2(_0581_),
    .B(_0583_),
    .C(_0584_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2727_ (.I(_2133_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2728_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[14].i3 ),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2729_ (.I(_0587_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2730_ (.A1(_0586_),
    .A2(_0567_),
    .B1(_0588_),
    .B2(_2207_),
    .C1(_2208_),
    .C2(_2366_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2731_ (.A1(_2258_),
    .A2(_0589_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2732_ (.A1(_2258_),
    .A2(_0585_),
    .B(_0590_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2733_ (.I(_0591_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2734_ (.I(_0592_),
    .ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2735_ (.A1(_2132_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.Y_CY[14].i3 ),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2736_ (.A1(_0587_),
    .A2(_2372_),
    .B1(_0593_),
    .B2(_2374_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2737_ (.A1(_0587_),
    .A2(_2260_),
    .A3(_0594_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2738_ (.I(_0595_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2739_ (.A1(_0587_),
    .A2(_2260_),
    .B(_0594_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2740_ (.A1(_0596_),
    .A2(_0597_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2741_ (.A1(_0578_),
    .A2(_0583_),
    .A3(_0584_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2742_ (.A1(_0598_),
    .A2(_0599_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2743_ (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[0].i2 ),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2744_ (.A1(_0586_),
    .A2(_0588_),
    .B1(_0601_),
    .B2(_2207_),
    .C1(_2208_),
    .C2(_0567_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2745_ (.I0(_0600_),
    .I1(_0602_),
    .S(_2248_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2746_ (.I(_0603_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2747_ (.I(_0604_),
    .ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2748_ (.A1(_0577_),
    .A2(_0598_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2749_ (.A1(_0562_),
    .A2(_0563_),
    .B(_0582_),
    .C(_0598_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2750_ (.A1(_0584_),
    .A2(_0596_),
    .A3(_0605_),
    .A4(_0606_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2751_ (.A1(\Arithmetic_Logic_Unit.ALU_001.Y_CY[0].i2 ),
    .A2(_2261_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2752_ (.A1(_2132_),
    .A2(_0601_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2753_ (.A1(_0601_),
    .A2(_2372_),
    .B1(_0609_),
    .B2(_2374_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2754_ (.A1(_0607_),
    .A2(_0608_),
    .A3(_0610_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2755_ (.I(_0601_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _2756_ (.A1(_0586_),
    .A2(_0612_),
    .B1(_2207_),
    .B2(_2118_),
    .C1(_2253_),
    .C2(_0588_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2757_ (.I0(_0611_),
    .I1(_0613_),
    .S(_2248_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2758_ (.I(_0614_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2759_ (.I(_0615_),
    .ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2760_ (.I(\Control_unit2.instr_decoder2.A[1] ),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2761_ (.A1(_2141_),
    .A2(\Arithmetic_Logic_Unit.ALU_001.p_Z ),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2762_ (.A1(\Control_unit2.instr_decoder2.A[2] ),
    .A2(_0617_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2763_ (.A1(_0616_),
    .A2(_0618_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2764_ (.I(_0619_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2765_ (.I(_0620_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2766_ (.I(_0620_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2767_ (.A1(\Control_unit1.instr_decoder1.A[0] ),
    .A2(\Control_unit1.instr_stage1[2] ),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2768_ (.A1(\Control_unit1.instr_stage1[1] ),
    .A2(_2115_),
    .A3(_0623_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2769_ (.A1(\Control_unit1.instr_stage1[0] ),
    .A2(_0624_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2770_ (.A1(\Control_unit1.instr_stage1[12] ),
    .A2(\Control_unit1.instr_stage1[11] ),
    .A3(_0625_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2771_ (.A1(\Control_unit1.instr_decoder1.A[2] ),
    .A2(\Control_unit1.instr_decoder1.A[1] ),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2772_ (.A1(_0626_),
    .A2(_0627_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2773_ (.A1(\Stack_pointer.SP[0] ),
    .A2(_0622_),
    .A3(_0628_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2774_ (.I(_0626_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2775_ (.I(_0627_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2776_ (.I(_0619_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2777_ (.A1(\Stack_pointer.SP[0] ),
    .A2(_0632_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2778_ (.A1(\Control_unit1.instr_stage1[3] ),
    .A2(_0630_),
    .B1(_0631_),
    .B2(_0633_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2779_ (.A1(\Stack_pointer.SP[0] ),
    .A2(_0621_),
    .B(_0629_),
    .C(_0634_),
    .ZN(\Stack_pointer.SP_next[0] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2780_ (.I(_0628_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2781_ (.A1(\Stack_pointer.SP[1] ),
    .A2(_0621_),
    .A3(_0635_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2782_ (.I(_0626_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2783_ (.I(_0637_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2784_ (.I(_0627_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2785_ (.I(_0639_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2786_ (.A1(\Stack_pointer.SP[1] ),
    .A2(_0622_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2787_ (.I(_0620_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2788_ (.A1(\Stack_pointer.SP[1] ),
    .A2(_0642_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2789_ (.A1(\Control_unit1.instr_stage1[4] ),
    .A2(_0638_),
    .B1(_0640_),
    .B2(_0641_),
    .C(_0643_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2790_ (.A1(_0636_),
    .A2(_0644_),
    .ZN(\Stack_pointer.SP_next[1] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2791_ (.A1(\Stack_pointer.SP[2] ),
    .A2(_0621_),
    .A3(_0635_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2792_ (.A1(\Stack_pointer.SP[2] ),
    .A2(_0622_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2793_ (.A1(\Stack_pointer.SP[2] ),
    .A2(_0642_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2794_ (.A1(\Control_unit1.instr_stage1[5] ),
    .A2(_0630_),
    .B1(_0631_),
    .B2(_0646_),
    .C(_0647_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2795_ (.A1(_0645_),
    .A2(_0648_),
    .ZN(\Stack_pointer.SP_next[2] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2796_ (.A1(\Stack_pointer.SP[3] ),
    .A2(_0621_),
    .A3(_0635_),
    .ZN(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2797_ (.A1(\Stack_pointer.SP[3] ),
    .A2(_0642_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2798_ (.I(_0619_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2799_ (.A1(\Stack_pointer.SP[3] ),
    .A2(_0651_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2800_ (.A1(\Control_unit1.instr_stage1[6] ),
    .A2(_0630_),
    .B1(_0631_),
    .B2(_0650_),
    .C(_0652_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2801_ (.A1(_0649_),
    .A2(_0653_),
    .ZN(\Stack_pointer.SP_next[3] ));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2802_ (.A1(\Stack_pointer.SP[4] ),
    .A2(_0622_),
    .A3(_0635_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2803_ (.A1(\Stack_pointer.SP[4] ),
    .A2(_0642_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2804_ (.A1(\Stack_pointer.SP[4] ),
    .A2(_0651_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2805_ (.A1(\Control_unit1.instr_stage1[7] ),
    .A2(_0630_),
    .B1(_0631_),
    .B2(_0655_),
    .C(_0656_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2806_ (.A1(_0654_),
    .A2(_0657_),
    .ZN(\Stack_pointer.SP_next[4] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2807_ (.A1(\Stack_pointer.SP[5] ),
    .A2(_0632_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2808_ (.A1(\Stack_pointer.SP[5] ),
    .A2(_0651_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2809_ (.A1(\Control_unit1.instr_stage1[8] ),
    .A2(_0637_),
    .B1(_0639_),
    .B2(_0658_),
    .C(_0659_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2810_ (.A1(_0638_),
    .A2(_0640_),
    .A3(_0658_),
    .B(_0660_),
    .ZN(\Stack_pointer.SP_next[5] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2811_ (.A1(\Stack_pointer.SP[6] ),
    .A2(_0632_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2812_ (.A1(\Stack_pointer.SP[6] ),
    .A2(_0651_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2813_ (.A1(\Control_unit1.instr_stage1[9] ),
    .A2(_0637_),
    .B1(_0639_),
    .B2(_0661_),
    .C(_0662_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2814_ (.A1(_0638_),
    .A2(_0640_),
    .A3(_0661_),
    .B(_0663_),
    .ZN(\Stack_pointer.SP_next[6] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2815_ (.A1(\Stack_pointer.SP[7] ),
    .A2(_0620_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2816_ (.A1(\Stack_pointer.SP[7] ),
    .A2(_0632_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2817_ (.A1(\Control_unit1.instr_stage1[10] ),
    .A2(_0637_),
    .B1(_0639_),
    .B2(_0664_),
    .C(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2818_ (.A1(_0638_),
    .A2(_0640_),
    .A3(_0664_),
    .B(_0666_),
    .ZN(\Stack_pointer.SP_next[7] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2819_ (.I(_0618_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2820_ (.A1(_2086_),
    .A2(_0667_),
    .B(_0616_),
    .ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2821_ (.I(\Control_unit1.instr_decoder1.A[2] ),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2822_ (.A1(_0668_),
    .A2(\Control_unit1.instr_decoder1.A[1] ),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2823_ (.A1(\Control_unit1.instr_decoder1.A[0] ),
    .A2(_0669_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2824_ (.I(_0670_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2825_ (.I(\Stack_pointer.SP[0] ),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2826_ (.A1(\Control_unit1.instr_stage1[12] ),
    .A2(\Control_unit1.instr_stage1[11] ),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2827_ (.A1(_0625_),
    .A2(_0673_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2828_ (.A1(_0672_),
    .A2(_0674_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2829_ (.A1(_0671_),
    .A2(_0675_),
    .B(\Control_unit1.instr_stage1[0] ),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2830_ (.A1(_0616_),
    .A2(_2086_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2831_ (.I(_0677_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2832_ (.A1(_2079_),
    .A2(_0678_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2833_ (.A1(_0633_),
    .A2(_0676_),
    .A3(_0679_),
    .ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2834_ (.I(_0677_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2835_ (.A1(_2084_),
    .A2(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2836_ (.I(_0670_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2837_ (.I(_0618_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2838_ (.A1(_0616_),
    .A2(_0683_),
    .B(_0674_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2839_ (.I(_0684_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2840_ (.A1(\Control_unit1.instr_stage1[1] ),
    .A2(_0682_),
    .B1(_0685_),
    .B2(\Stack_pointer.SP[1] ),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2841_ (.A1(_0681_),
    .A2(_0686_),
    .ZN(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2842_ (.I(_2101_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2843_ (.I(_0687_),
    .Z(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _2844_ (.A1(_0688_),
    .A2(_0678_),
    .B1(_0671_),
    .B2(\Control_unit1.instr_stage1[2] ),
    .C1(_0684_),
    .C2(\Stack_pointer.SP[2] ),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2845_ (.I(_0689_),
    .ZN(net40));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2846_ (.A1(\Control_unit2.instr_stage2[3] ),
    .A2(_0680_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2847_ (.A1(\Control_unit1.instr_stage1[3] ),
    .A2(_0682_),
    .B1(_0685_),
    .B2(\Stack_pointer.SP[3] ),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2848_ (.A1(_0690_),
    .A2(_0691_),
    .ZN(net41));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2849_ (.A1(\Control_unit2.instr_stage2[4] ),
    .A2(_0680_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2850_ (.A1(\Control_unit1.instr_stage1[4] ),
    .A2(_0682_),
    .B1(_0685_),
    .B2(\Stack_pointer.SP[4] ),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2851_ (.A1(_0692_),
    .A2(_0693_),
    .ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2852_ (.A1(\Control_unit2.instr_stage2[5] ),
    .A2(_0680_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2853_ (.A1(\Control_unit1.instr_stage1[5] ),
    .A2(_0682_),
    .B1(_0685_),
    .B2(\Stack_pointer.SP[5] ),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2854_ (.A1(_0694_),
    .A2(_0695_),
    .ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2855_ (.A1(\Control_unit2.instr_stage2[6] ),
    .A2(_0678_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2856_ (.A1(\Control_unit1.instr_stage1[6] ),
    .A2(_0671_),
    .B1(_0684_),
    .B2(\Stack_pointer.SP[6] ),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2857_ (.A1(_0696_),
    .A2(_0697_),
    .ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2858_ (.A1(\Control_unit2.instr_stage2[7] ),
    .A2(_0678_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2859_ (.A1(\Control_unit1.instr_stage1[7] ),
    .A2(_0671_),
    .B1(_0684_),
    .B2(\Stack_pointer.SP[7] ),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2860_ (.A1(_0698_),
    .A2(_0699_),
    .ZN(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2861_ (.I(\Control_unit2.instr_stage2[12] ),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2862_ (.I(\Arithmetic_Logic_Unit.ALU_001.p_Z ),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2863_ (.A1(_0700_),
    .A2(\Control_unit2.instr_stage2[11] ),
    .B(_0701_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2864_ (.I(\Control_unit2.instr_stage2[11] ),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2865_ (.A1(_2089_),
    .A2(_0703_),
    .B(\Arithmetic_Logic_Unit.ALU_001.p_Z ),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2866_ (.A1(_2088_),
    .A2(_0702_),
    .A3(_0704_),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2867_ (.I(_0705_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2868_ (.A1(net70),
    .A2(_0706_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2869_ (.A1(_2088_),
    .A2(_2090_),
    .B(net35),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2870_ (.I(_0708_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2871_ (.I(_0709_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2872_ (.I(_0683_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2873_ (.I(_0711_),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2874_ (.A1(_0683_),
    .A2(_0705_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2875_ (.I(_0713_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2876_ (.A1(net47),
    .A2(net51),
    .A3(net52),
    .A4(net53),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2877_ (.A1(net54),
    .A2(_0715_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2878_ (.A1(\Control_unit2.instr_stage2[4] ),
    .A2(_0712_),
    .B1(_0714_),
    .B2(_0716_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2879_ (.A1(net35),
    .A2(net46),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2880_ (.I(_0718_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2881_ (.I(net54),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2882_ (.A1(_0707_),
    .A2(_0710_),
    .A3(_0717_),
    .B1(_0719_),
    .B2(_0720_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2883_ (.I(_0709_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2884_ (.A1(net54),
    .A2(_0715_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2885_ (.A1(net55),
    .A2(_0722_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2886_ (.A1(net55),
    .A2(_0722_),
    .Z(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2887_ (.A1(_0723_),
    .A2(_0724_),
    .B(_0714_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2888_ (.I(_0705_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2889_ (.A1(\Control_unit2.instr_stage2[5] ),
    .A2(_0712_),
    .B1(_0726_),
    .B2(_2274_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2890_ (.I(net55),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2891_ (.A1(_0721_),
    .A2(_0725_),
    .A3(_0727_),
    .B1(_0719_),
    .B2(_0728_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2892_ (.I(net56),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2893_ (.I(_0718_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2894_ (.A1(_0683_),
    .A2(_0705_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2895_ (.I(_0731_),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2896_ (.A1(net56),
    .A2(_0723_),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2897_ (.A1(_0732_),
    .A2(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2898_ (.A1(\Control_unit2.instr_stage2[6] ),
    .A2(_0712_),
    .B1(_0706_),
    .B2(_2250_),
    .C(_0734_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2899_ (.A1(_0729_),
    .A2(_0730_),
    .B1(_0710_),
    .B2(_0735_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2900_ (.I(net57),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2901_ (.A1(net55),
    .A2(net56),
    .A3(_0722_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2902_ (.A1(net57),
    .A2(_0737_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2903_ (.A1(_0731_),
    .A2(_0738_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2904_ (.A1(\Control_unit2.instr_stage2[7] ),
    .A2(_0712_),
    .B1(_0706_),
    .B2(_2273_),
    .C(_0739_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2905_ (.A1(_0736_),
    .A2(_0719_),
    .B1(_0710_),
    .B2(_0740_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2906_ (.A1(_0736_),
    .A2(_0737_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2907_ (.A1(net58),
    .A2(_0741_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2908_ (.I(net58),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2909_ (.A1(_0736_),
    .A2(_0737_),
    .B(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2910_ (.A1(_0742_),
    .A2(_0744_),
    .B(_0714_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2911_ (.I(\Control_unit2.instr_stage2[8] ),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2912_ (.I(_0711_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2913_ (.A1(_0746_),
    .A2(_0747_),
    .B1(_0726_),
    .B2(_2283_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2914_ (.I(_0718_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2915_ (.A1(_0721_),
    .A2(_0745_),
    .A3(_0748_),
    .B1(_0749_),
    .B2(_0743_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2916_ (.I(net59),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2917_ (.I(\Control_unit2.instr_stage2[9] ),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2918_ (.A1(_2088_),
    .A2(_0702_),
    .A3(_0704_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2919_ (.I(_0752_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2920_ (.A1(net59),
    .A2(_0742_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2921_ (.A1(_2335_),
    .A2(_0753_),
    .B1(_0732_),
    .B2(_0754_),
    .C(_0709_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2922_ (.A1(_0751_),
    .A2(_0667_),
    .B(_0755_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2923_ (.A1(_0750_),
    .A2(_0730_),
    .B(_0756_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2924_ (.A1(_2341_),
    .A2(_2353_),
    .B(_0726_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2925_ (.I(\Control_unit2.instr_stage2[10] ),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2926_ (.I(net48),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2927_ (.A1(net58),
    .A2(net59),
    .A3(_0741_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2928_ (.A1(_0759_),
    .A2(_0760_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2929_ (.A1(_0758_),
    .A2(_0747_),
    .B1(_0714_),
    .B2(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2930_ (.A1(_0721_),
    .A2(_0757_),
    .A3(_0762_),
    .B1(_0749_),
    .B2(_0759_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2931_ (.A1(net62),
    .A2(_0706_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2932_ (.I(\Control_unit2.instr_stage2[11] ),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2933_ (.A1(_0759_),
    .A2(_0760_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2934_ (.A1(net49),
    .A2(_0765_),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2935_ (.A1(_0764_),
    .A2(_0747_),
    .B1(_0713_),
    .B2(_0766_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2936_ (.I(net49),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2937_ (.A1(_0721_),
    .A2(_0763_),
    .A3(_0767_),
    .B1(_0749_),
    .B2(_0768_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2938_ (.I(net50),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2939_ (.A1(net49),
    .A2(_0765_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2940_ (.A1(net50),
    .A2(_0770_),
    .Z(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2941_ (.A1(_0711_),
    .A2(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2942_ (.A1(_2089_),
    .A2(_0711_),
    .B(_0772_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2943_ (.I0(_0571_),
    .I1(_0773_),
    .S(_0726_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2944_ (.A1(_0769_),
    .A2(_0719_),
    .B1(_0710_),
    .B2(_0774_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2945_ (.A1(\Control_unit1.instr_stage1[0] ),
    .A2(_0673_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2946_ (.A1(_0624_),
    .A2(_0775_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2947_ (.A1(_0669_),
    .A2(_0776_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2948_ (.I(_0777_),
    .Z(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2949_ (.I(_0778_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2950_ (.I(net18),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2951_ (.I(_0780_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2952_ (.I(_0777_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2953_ (.I(_0782_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2954_ (.A1(_0781_),
    .A2(_0783_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2955_ (.A1(_2146_),
    .A2(_0779_),
    .B(_0784_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2956_ (.I(net25),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2957_ (.I(_0785_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2958_ (.A1(_0786_),
    .A2(_0783_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2959_ (.A1(_2172_),
    .A2(_0779_),
    .B(_0787_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2960_ (.I(net26),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2961_ (.I(_0788_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2962_ (.A1(_0789_),
    .A2(_0783_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2963_ (.A1(_2190_),
    .A2(_0779_),
    .B(_0790_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2964_ (.I(net27),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2965_ (.I(_0791_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2966_ (.A1(_0792_),
    .A2(_0783_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2967_ (.A1(_2212_),
    .A2(_0779_),
    .B(_0793_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2968_ (.I(_2232_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2969_ (.I(_0794_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2970_ (.I(_0778_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2971_ (.I(net28),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2972_ (.I(_0797_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2973_ (.I(_0782_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2974_ (.A1(_0798_),
    .A2(_0799_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2975_ (.A1(_0795_),
    .A2(_0796_),
    .B(_0800_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2976_ (.I(net29),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2977_ (.I(_0801_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2978_ (.A1(_0802_),
    .A2(_0799_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2979_ (.A1(_2257_),
    .A2(_0796_),
    .B(_0803_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2980_ (.I(net30),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2981_ (.I(_0804_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2982_ (.A1(_0805_),
    .A2(_0799_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2983_ (.A1(_2278_),
    .A2(_0796_),
    .B(_0806_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2984_ (.I(net31),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2985_ (.I(_0807_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2986_ (.A1(_0808_),
    .A2(_0799_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2987_ (.A1(_2298_),
    .A2(_0796_),
    .B(_0809_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2988_ (.I(_0778_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2989_ (.I(net32),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2990_ (.I(_0811_),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2991_ (.I(_0782_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2992_ (.A1(_0812_),
    .A2(_0813_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2993_ (.A1(_2322_),
    .A2(_0810_),
    .B(_0814_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2994_ (.I(net33),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2995_ (.I(_0815_),
    .Z(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2996_ (.A1(_0816_),
    .A2(_0813_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2997_ (.A1(_2336_),
    .A2(_0810_),
    .B(_0817_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2998_ (.I(net19),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2999_ (.I(_0818_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3000_ (.A1(_0819_),
    .A2(_0813_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3001_ (.A1(_2355_),
    .A2(_0810_),
    .B(_0820_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3002_ (.I(_2370_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3003_ (.I(_0821_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3004_ (.I(net20),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3005_ (.I(_0823_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3006_ (.A1(_0824_),
    .A2(_0813_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3007_ (.A1(_0822_),
    .A2(_0810_),
    .B(_0825_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3008_ (.I(_0778_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3009_ (.I(net21),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3010_ (.I(_0827_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3011_ (.I(_0782_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3012_ (.A1(_0828_),
    .A2(_0829_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3013_ (.A1(_0572_),
    .A2(_0826_),
    .B(_0830_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3014_ (.I(net22),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3015_ (.I(_0831_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3016_ (.A1(_0832_),
    .A2(_0829_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3017_ (.A1(_0592_),
    .A2(_0826_),
    .B(_0833_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3018_ (.I(net23),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3019_ (.I(_0834_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3020_ (.A1(_0835_),
    .A2(_0829_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3021_ (.A1(_0604_),
    .A2(_0826_),
    .B(_0836_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3022_ (.I(net24),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3023_ (.I(_0837_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3024_ (.A1(_0838_),
    .A2(_0829_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3025_ (.A1(_0615_),
    .A2(_0826_),
    .B(_0839_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3026_ (.A1(\Control_unit1.instr_decoder1.A[2] ),
    .A2(\Control_unit1.instr_decoder1.A[1] ),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3027_ (.A1(_0840_),
    .A2(_0623_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3028_ (.I(_0841_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3029_ (.I(_0842_),
    .Z(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3030_ (.I(_0841_),
    .Z(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3031_ (.A1(_0780_),
    .A2(_0844_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3032_ (.A1(_2097_),
    .A2(_0843_),
    .B(_0845_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3033_ (.A1(_0785_),
    .A2(_0844_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3034_ (.A1(_2151_),
    .A2(_0843_),
    .B(_0846_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3035_ (.A1(_0788_),
    .A2(_0844_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3036_ (.A1(_2177_),
    .A2(_0843_),
    .B(_0847_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3037_ (.I(_0841_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3038_ (.A1(_0791_),
    .A2(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3039_ (.A1(_2193_),
    .A2(_0843_),
    .B(_0849_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3040_ (.I0(_0798_),
    .I1(_2206_),
    .S(_0848_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3041_ (.I(_0850_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3042_ (.I0(_0802_),
    .I1(_2274_),
    .S(_0848_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3043_ (.I(_0851_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3044_ (.I(_0842_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3045_ (.I0(_0805_),
    .I1(_2250_),
    .S(_0852_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3046_ (.I(_0853_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3047_ (.I0(_0808_),
    .I1(_2273_),
    .S(_0852_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3048_ (.I(_0854_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3049_ (.I0(_0812_),
    .I1(_2283_),
    .S(_0852_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3050_ (.I(_0855_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3051_ (.I0(_0816_),
    .I1(_2318_),
    .S(_0852_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3052_ (.I(_0856_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3053_ (.A1(_0818_),
    .A2(_0848_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3054_ (.A1(_2338_),
    .A2(_0844_),
    .B(_0857_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3055_ (.I(_0842_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3056_ (.I0(_0824_),
    .I1(_2337_),
    .S(_0858_),
    .Z(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3057_ (.I(_0859_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3058_ (.I0(_0828_),
    .I1(_2366_),
    .S(_0858_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3059_ (.I(_0860_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3060_ (.I0(_0832_),
    .I1(_0567_),
    .S(_0858_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3061_ (.I(_0861_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3062_ (.I0(_0835_),
    .I1(_0588_),
    .S(_0858_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3063_ (.I(_0862_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3064_ (.I0(_0838_),
    .I1(_0612_),
    .S(_0842_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3065_ (.I(_0863_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3066_ (.A1(_0687_),
    .A2(_2233_),
    .B(\Control_unit2.instr_decoder2.A[2] ),
    .C(\Control_unit2.instr_decoder2.A[1] ),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3067_ (.I(_2233_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3068_ (.A1(_2106_),
    .A2(_2251_),
    .B1(_2253_),
    .B2(_0612_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3069_ (.A1(_0865_),
    .A2(_0866_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3070_ (.A1(_0864_),
    .A2(_0867_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3071_ (.I(_0610_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3072_ (.A1(_0608_),
    .A2(_0869_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3073_ (.A1(_0596_),
    .A2(_0606_),
    .B(_0870_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3074_ (.A1(_0584_),
    .A2(_0605_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3075_ (.A1(_0612_),
    .A2(_2261_),
    .A3(_0610_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3076_ (.A1(_0872_),
    .A2(_0873_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3077_ (.A1(_0871_),
    .A2(_0874_),
    .B(_0688_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3078_ (.A1(_0688_),
    .A2(_0871_),
    .A3(_0874_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3079_ (.A1(_0865_),
    .A2(_0875_),
    .A3(_0876_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3080_ (.A1(_2121_),
    .A2(_0864_),
    .B1(_0868_),
    .B2(_0877_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3081_ (.A1(\Control_unit2.instr_stage2[9] ),
    .A2(\Control_unit2.instr_stage2[10] ),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3082_ (.A1(_0746_),
    .A2(_0878_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3083_ (.A1(_0687_),
    .A2(\Control_unit2.instr_decoder2.A[1] ),
    .B(_2141_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3084_ (.A1(_2119_),
    .A2(_2087_),
    .B1(_0880_),
    .B2(_2085_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3085_ (.A1(_0700_),
    .A2(_0764_),
    .A3(_0881_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3086_ (.I(_0882_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3087_ (.A1(_0879_),
    .A2(_0883_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3088_ (.I(_0884_),
    .Z(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3089_ (.I(_0885_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3090_ (.I(_0884_),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3091_ (.I(_0887_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3092_ (.A1(_0781_),
    .A2(_0888_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3093_ (.A1(_2146_),
    .A2(_0886_),
    .B(_0889_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3094_ (.A1(_0786_),
    .A2(_0888_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3095_ (.A1(_2172_),
    .A2(_0886_),
    .B(_0890_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3096_ (.A1(_0789_),
    .A2(_0888_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3097_ (.A1(_2190_),
    .A2(_0886_),
    .B(_0891_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3098_ (.A1(_0792_),
    .A2(_0888_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3099_ (.A1(_2212_),
    .A2(_0886_),
    .B(_0892_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3100_ (.I(_0885_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3101_ (.I(_0887_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3102_ (.A1(_0798_),
    .A2(_0894_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3103_ (.A1(_0795_),
    .A2(_0893_),
    .B(_0895_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3104_ (.A1(_0802_),
    .A2(_0894_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3105_ (.A1(_2257_),
    .A2(_0893_),
    .B(_0896_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3106_ (.A1(_0805_),
    .A2(_0894_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3107_ (.A1(_2278_),
    .A2(_0893_),
    .B(_0897_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3108_ (.A1(_0808_),
    .A2(_0894_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3109_ (.A1(_2298_),
    .A2(_0893_),
    .B(_0898_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3110_ (.I(_0885_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3111_ (.I(_0887_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3112_ (.A1(_0812_),
    .A2(_0900_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3113_ (.A1(_2322_),
    .A2(_0899_),
    .B(_0901_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3114_ (.A1(_0816_),
    .A2(_0900_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3115_ (.A1(_2336_),
    .A2(_0899_),
    .B(_0902_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3116_ (.A1(_0819_),
    .A2(_0900_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3117_ (.A1(_2355_),
    .A2(_0899_),
    .B(_0903_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3118_ (.A1(_0824_),
    .A2(_0900_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3119_ (.A1(_0822_),
    .A2(_0899_),
    .B(_0904_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3120_ (.I(_0885_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3121_ (.I(_0887_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3122_ (.A1(_0828_),
    .A2(_0906_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3123_ (.A1(_0572_),
    .A2(_0905_),
    .B(_0907_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3124_ (.A1(_0832_),
    .A2(_0906_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3125_ (.A1(_0592_),
    .A2(_0905_),
    .B(_0908_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3126_ (.A1(_0835_),
    .A2(_0906_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3127_ (.A1(_0604_),
    .A2(_0905_),
    .B(_0909_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3128_ (.A1(_0838_),
    .A2(_0906_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3129_ (.A1(_0615_),
    .A2(_0905_),
    .B(_0910_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3130_ (.A1(_2349_),
    .A2(_2352_),
    .B1(_0561_),
    .B2(_0564_),
    .C(_2332_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3131_ (.A1(_2312_),
    .A2(_2313_),
    .B(_2314_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3132_ (.A1(_2300_),
    .A2(_2303_),
    .A3(_2309_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3133_ (.A1(_2241_),
    .A2(_2246_),
    .B1(_2269_),
    .B2(_2270_),
    .C1(_0912_),
    .C2(_0913_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3134_ (.A1(_0687_),
    .A2(_2251_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3135_ (.A1(_2129_),
    .A2(_0915_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3136_ (.A1(_2161_),
    .A2(_2183_),
    .A3(_2228_),
    .A4(_0916_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3137_ (.A1(_2204_),
    .A2(_2295_),
    .A3(_0914_),
    .A4(_0917_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3138_ (.A1(_2364_),
    .A2(_0585_),
    .A3(_0911_),
    .A4(_0918_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3139_ (.A1(_0600_),
    .A2(_0919_),
    .B(_0865_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3140_ (.A1(_2206_),
    .A2(_2274_),
    .A3(_2250_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3141_ (.A1(_2084_),
    .A2(_2135_),
    .A3(_2165_),
    .A4(_2185_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3142_ (.A1(_0921_),
    .A2(_0922_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3143_ (.A1(_2319_),
    .A2(_2333_),
    .A3(_2340_),
    .A4(_2368_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3144_ (.A1(_2285_),
    .A2(_0923_),
    .A3(_0924_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3145_ (.A1(_0568_),
    .A2(_0589_),
    .A3(_0602_),
    .A4(_0925_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3146_ (.A1(_2140_),
    .A2(_0613_),
    .A3(_0926_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3147_ (.A1(_0586_),
    .A2(_0701_),
    .B(_0927_),
    .C(_2233_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3148_ (.A1(_0865_),
    .A2(_0611_),
    .B(_0864_),
    .C(_0928_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3149_ (.A1(_0701_),
    .A2(_0864_),
    .B1(_0920_),
    .B2(_0929_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3150_ (.I(\Control_unit2.instr_stage2[8] ),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3151_ (.A1(_0930_),
    .A2(\Control_unit2.instr_stage2[9] ),
    .A3(\Control_unit2.instr_stage2[10] ),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3152_ (.A1(_2089_),
    .A2(_0764_),
    .A3(_0881_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3153_ (.I(_0932_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3154_ (.A1(_0931_),
    .A2(_0933_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3155_ (.I(_0934_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3156_ (.I(_0935_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3157_ (.I(_0934_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3158_ (.I(_0937_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3159_ (.A1(_0781_),
    .A2(_0938_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3160_ (.A1(_2146_),
    .A2(_0936_),
    .B(_0939_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3161_ (.A1(_0786_),
    .A2(_0938_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3162_ (.A1(_2172_),
    .A2(_0936_),
    .B(_0940_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3163_ (.A1(_0789_),
    .A2(_0938_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3164_ (.A1(_2190_),
    .A2(_0936_),
    .B(_0941_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3165_ (.A1(_0792_),
    .A2(_0938_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3166_ (.A1(_2212_),
    .A2(_0936_),
    .B(_0942_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3167_ (.I(_0935_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3168_ (.I(_0937_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3169_ (.A1(_0798_),
    .A2(_0944_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3170_ (.A1(_0795_),
    .A2(_0943_),
    .B(_0945_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3171_ (.A1(_0802_),
    .A2(_0944_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3172_ (.A1(_2257_),
    .A2(_0943_),
    .B(_0946_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3173_ (.A1(_0805_),
    .A2(_0944_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3174_ (.A1(_2278_),
    .A2(_0943_),
    .B(_0947_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3175_ (.A1(_0808_),
    .A2(_0944_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3176_ (.A1(_2298_),
    .A2(_0943_),
    .B(_0948_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3177_ (.I(_0935_),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3178_ (.I(_0937_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3179_ (.A1(_0812_),
    .A2(_0950_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3180_ (.A1(_2322_),
    .A2(_0949_),
    .B(_0951_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3181_ (.A1(_0816_),
    .A2(_0950_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3182_ (.A1(_2336_),
    .A2(_0949_),
    .B(_0952_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3183_ (.A1(_0819_),
    .A2(_0950_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3184_ (.A1(_2355_),
    .A2(_0949_),
    .B(_0953_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3185_ (.A1(_0824_),
    .A2(_0950_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3186_ (.A1(_0822_),
    .A2(_0949_),
    .B(_0954_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3187_ (.I(_0935_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3188_ (.I(_0937_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3189_ (.A1(_0828_),
    .A2(_0956_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3190_ (.A1(_0572_),
    .A2(_0955_),
    .B(_0957_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3191_ (.A1(_0832_),
    .A2(_0956_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3192_ (.A1(_0592_),
    .A2(_0955_),
    .B(_0958_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3193_ (.A1(_0835_),
    .A2(_0956_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3194_ (.A1(_0604_),
    .A2(_0955_),
    .B(_0959_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3195_ (.A1(_0838_),
    .A2(_0956_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3196_ (.A1(_0615_),
    .A2(_0955_),
    .B(_0960_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3197_ (.I(_2145_),
    .Z(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3198_ (.I(_0961_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3199_ (.I(\Control_unit2.instr_stage2[10] ),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3200_ (.A1(_0930_),
    .A2(_0751_),
    .A3(_0963_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3201_ (.A1(_2090_),
    .A2(_0881_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3202_ (.I(_0965_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3203_ (.A1(_0964_),
    .A2(_0966_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3204_ (.I(_0967_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3205_ (.I(_0968_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3206_ (.I(_0967_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3207_ (.I(_0970_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3208_ (.A1(_0781_),
    .A2(_0971_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3209_ (.A1(_0962_),
    .A2(_0969_),
    .B(_0972_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3210_ (.I(_2171_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3211_ (.I(_0973_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3212_ (.A1(_0786_),
    .A2(_0971_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3213_ (.A1(_0974_),
    .A2(_0969_),
    .B(_0975_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3214_ (.I(_2189_),
    .Z(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3215_ (.I(_0976_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3216_ (.A1(_0789_),
    .A2(_0971_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3217_ (.A1(_0977_),
    .A2(_0969_),
    .B(_0978_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3218_ (.I(_2211_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3219_ (.I(_0979_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3220_ (.A1(_0792_),
    .A2(_0971_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3221_ (.A1(_0980_),
    .A2(_0969_),
    .B(_0981_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3222_ (.I(_0968_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3223_ (.I(_0797_),
    .Z(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3224_ (.I(_0970_),
    .Z(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3225_ (.A1(_0983_),
    .A2(_0984_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3226_ (.A1(_0795_),
    .A2(_0982_),
    .B(_0985_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3227_ (.I(_2256_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3228_ (.I(_0986_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3229_ (.I(_0801_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3230_ (.A1(_0988_),
    .A2(_0984_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3231_ (.A1(_0987_),
    .A2(_0982_),
    .B(_0989_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3232_ (.I(_2277_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3233_ (.I(_0990_),
    .Z(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3234_ (.I(_0804_),
    .Z(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3235_ (.A1(_0992_),
    .A2(_0984_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3236_ (.A1(_0991_),
    .A2(_0982_),
    .B(_0993_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3237_ (.I(_2297_),
    .Z(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3238_ (.I(_0994_),
    .Z(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3239_ (.I(_0807_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3240_ (.A1(_0996_),
    .A2(_0984_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3241_ (.A1(_0995_),
    .A2(_0982_),
    .B(_0997_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3242_ (.I(_2321_),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3243_ (.I(_0998_),
    .Z(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3244_ (.I(_0968_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3245_ (.I(_0811_),
    .Z(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3246_ (.I(_0970_),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3247_ (.A1(_1001_),
    .A2(_1002_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3248_ (.A1(_0999_),
    .A2(_1000_),
    .B(_1003_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3249_ (.I(_2335_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3250_ (.I(_1004_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3251_ (.I(_0815_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3252_ (.A1(_1006_),
    .A2(_1002_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3253_ (.A1(_1005_),
    .A2(_1000_),
    .B(_1007_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3254_ (.I(_2354_),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3255_ (.I(_1008_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3256_ (.A1(_0819_),
    .A2(_1002_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3257_ (.A1(_1009_),
    .A2(_1000_),
    .B(_1010_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3258_ (.I(_0823_),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3259_ (.A1(_1011_),
    .A2(_1002_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3260_ (.A1(_0822_),
    .A2(_1000_),
    .B(_1012_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3261_ (.I(_0571_),
    .Z(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3262_ (.I(_1013_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3263_ (.I(_0968_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3264_ (.I(_0827_),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3265_ (.I(_0970_),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3266_ (.A1(_1016_),
    .A2(_1017_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3267_ (.A1(_1014_),
    .A2(_1015_),
    .B(_1018_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3268_ (.I(_0591_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3269_ (.I(_1019_),
    .Z(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3270_ (.I(_0831_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3271_ (.A1(_1021_),
    .A2(_1017_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3272_ (.A1(_1020_),
    .A2(_1015_),
    .B(_1022_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3273_ (.I(_0603_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3274_ (.I(_1023_),
    .Z(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3275_ (.I(_0834_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3276_ (.A1(_1025_),
    .A2(_1017_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3277_ (.A1(_1024_),
    .A2(_1015_),
    .B(_1026_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3278_ (.I(_0614_),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3279_ (.I(_1027_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3280_ (.I(_0837_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3281_ (.A1(_1029_),
    .A2(_1017_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3282_ (.A1(_1028_),
    .A2(_1015_),
    .B(_1030_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3283_ (.I(_0932_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3284_ (.I(\Control_unit2.instr_stage2[9] ),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3285_ (.A1(_0930_),
    .A2(_1032_),
    .A3(_0758_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3286_ (.A1(_1031_),
    .A2(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3287_ (.I(_1034_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3288_ (.I(_1035_),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3289_ (.I(_0780_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3290_ (.I(_1034_),
    .Z(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3291_ (.I(_1038_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3292_ (.A1(_1037_),
    .A2(_1039_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3293_ (.A1(_0962_),
    .A2(_1036_),
    .B(_1040_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3294_ (.I(_0785_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3295_ (.A1(_1041_),
    .A2(_1039_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3296_ (.A1(_0974_),
    .A2(_1036_),
    .B(_1042_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3297_ (.I(_0788_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3298_ (.A1(_1043_),
    .A2(_1039_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3299_ (.A1(_0977_),
    .A2(_1036_),
    .B(_1044_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3300_ (.I(_0791_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3301_ (.A1(_1045_),
    .A2(_1039_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3302_ (.A1(_0980_),
    .A2(_1036_),
    .B(_1046_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3303_ (.I(_0794_),
    .Z(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3304_ (.I(_1035_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3305_ (.I(_1038_),
    .Z(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3306_ (.A1(_0983_),
    .A2(_1049_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3307_ (.A1(_1047_),
    .A2(_1048_),
    .B(_1050_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3308_ (.A1(_0988_),
    .A2(_1049_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3309_ (.A1(_0987_),
    .A2(_1048_),
    .B(_1051_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3310_ (.A1(_0992_),
    .A2(_1049_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3311_ (.A1(_0991_),
    .A2(_1048_),
    .B(_1052_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3312_ (.A1(_0996_),
    .A2(_1049_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3313_ (.A1(_0995_),
    .A2(_1048_),
    .B(_1053_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3314_ (.I(_1035_),
    .Z(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3315_ (.I(_1038_),
    .Z(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3316_ (.A1(_1001_),
    .A2(_1055_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3317_ (.A1(_0999_),
    .A2(_1054_),
    .B(_1056_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3318_ (.A1(_1006_),
    .A2(_1055_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3319_ (.A1(_1005_),
    .A2(_1054_),
    .B(_1057_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3320_ (.I(_0818_),
    .Z(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3321_ (.A1(_1058_),
    .A2(_1055_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3322_ (.A1(_1009_),
    .A2(_1054_),
    .B(_1059_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3323_ (.I(_0821_),
    .Z(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3324_ (.A1(_1011_),
    .A2(_1055_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3325_ (.A1(_1060_),
    .A2(_1054_),
    .B(_1061_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3326_ (.I(_1035_),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3327_ (.I(_1038_),
    .Z(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3328_ (.A1(_1016_),
    .A2(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3329_ (.A1(_1014_),
    .A2(_1062_),
    .B(_1064_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3330_ (.A1(_1021_),
    .A2(_1063_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3331_ (.A1(_1020_),
    .A2(_1062_),
    .B(_1065_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3332_ (.A1(_1025_),
    .A2(_1063_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3333_ (.A1(_1024_),
    .A2(_1062_),
    .B(_1066_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3334_ (.A1(_1029_),
    .A2(_1063_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3335_ (.A1(_1028_),
    .A2(_1062_),
    .B(_1067_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3336_ (.A1(_0746_),
    .A2(_0751_),
    .A3(_0963_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3337_ (.A1(_1031_),
    .A2(_1068_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3338_ (.I(_1069_),
    .Z(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3339_ (.I(_1070_),
    .Z(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3340_ (.I(_1069_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3341_ (.I(_1072_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3342_ (.A1(_1037_),
    .A2(_1073_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3343_ (.A1(_0962_),
    .A2(_1071_),
    .B(_1074_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3344_ (.A1(_1041_),
    .A2(_1073_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3345_ (.A1(_0974_),
    .A2(_1071_),
    .B(_1075_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3346_ (.A1(_1043_),
    .A2(_1073_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3347_ (.A1(_0977_),
    .A2(_1071_),
    .B(_1076_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3348_ (.A1(_1045_),
    .A2(_1073_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3349_ (.A1(_0980_),
    .A2(_1071_),
    .B(_1077_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3350_ (.I(_1070_),
    .Z(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3351_ (.I(_1072_),
    .Z(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3352_ (.A1(_0983_),
    .A2(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3353_ (.A1(_1047_),
    .A2(_1078_),
    .B(_1080_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3354_ (.A1(_0988_),
    .A2(_1079_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3355_ (.A1(_0987_),
    .A2(_1078_),
    .B(_1081_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3356_ (.A1(_0992_),
    .A2(_1079_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3357_ (.A1(_0991_),
    .A2(_1078_),
    .B(_1082_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3358_ (.A1(_0996_),
    .A2(_1079_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3359_ (.A1(_0995_),
    .A2(_1078_),
    .B(_1083_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3360_ (.I(_1070_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3361_ (.I(_1072_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3362_ (.A1(_1001_),
    .A2(_1085_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3363_ (.A1(_0999_),
    .A2(_1084_),
    .B(_1086_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3364_ (.A1(_1006_),
    .A2(_1085_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3365_ (.A1(_1005_),
    .A2(_1084_),
    .B(_1087_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3366_ (.A1(_1058_),
    .A2(_1085_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3367_ (.A1(_1009_),
    .A2(_1084_),
    .B(_1088_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3368_ (.A1(_1011_),
    .A2(_1085_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3369_ (.A1(_1060_),
    .A2(_1084_),
    .B(_1089_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3370_ (.I(_1070_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3371_ (.I(_1072_),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3372_ (.A1(_1016_),
    .A2(_1091_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3373_ (.A1(_1014_),
    .A2(_1090_),
    .B(_1092_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3374_ (.A1(_1021_),
    .A2(_1091_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3375_ (.A1(_1020_),
    .A2(_1090_),
    .B(_1093_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3376_ (.A1(_1025_),
    .A2(_1091_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3377_ (.A1(_1024_),
    .A2(_1090_),
    .B(_1094_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3378_ (.A1(_1029_),
    .A2(_1091_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3379_ (.A1(_1028_),
    .A2(_1090_),
    .B(_1095_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3380_ (.A1(_1031_),
    .A2(_0964_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3381_ (.I(_1096_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3382_ (.I(_1097_),
    .Z(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3383_ (.I(_1096_),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3384_ (.I(_1099_),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3385_ (.A1(_1037_),
    .A2(_1100_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3386_ (.A1(_0962_),
    .A2(_1098_),
    .B(_1101_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3387_ (.A1(_1041_),
    .A2(_1100_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3388_ (.A1(_0974_),
    .A2(_1098_),
    .B(_1102_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3389_ (.A1(_1043_),
    .A2(_1100_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3390_ (.A1(_0977_),
    .A2(_1098_),
    .B(_1103_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3391_ (.A1(_1045_),
    .A2(_1100_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3392_ (.A1(_0980_),
    .A2(_1098_),
    .B(_1104_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3393_ (.I(_1097_),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3394_ (.I(_1099_),
    .Z(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3395_ (.A1(_0983_),
    .A2(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3396_ (.A1(_1047_),
    .A2(_1105_),
    .B(_1107_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3397_ (.A1(_0988_),
    .A2(_1106_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3398_ (.A1(_0987_),
    .A2(_1105_),
    .B(_1108_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3399_ (.A1(_0992_),
    .A2(_1106_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3400_ (.A1(_0991_),
    .A2(_1105_),
    .B(_1109_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3401_ (.A1(_0996_),
    .A2(_1106_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3402_ (.A1(_0995_),
    .A2(_1105_),
    .B(_1110_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3403_ (.I(_1097_),
    .Z(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3404_ (.I(_1099_),
    .Z(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3405_ (.A1(_1001_),
    .A2(_1112_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3406_ (.A1(_0999_),
    .A2(_1111_),
    .B(_1113_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3407_ (.A1(_1006_),
    .A2(_1112_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3408_ (.A1(_1005_),
    .A2(_1111_),
    .B(_1114_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3409_ (.A1(_1058_),
    .A2(_1112_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3410_ (.A1(_1009_),
    .A2(_1111_),
    .B(_1115_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3411_ (.A1(_1011_),
    .A2(_1112_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3412_ (.A1(_1060_),
    .A2(_1111_),
    .B(_1116_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3413_ (.I(_1097_),
    .Z(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3414_ (.I(_1099_),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3415_ (.A1(_1016_),
    .A2(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3416_ (.A1(_1014_),
    .A2(_1117_),
    .B(_1119_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3417_ (.A1(_1021_),
    .A2(_1118_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3418_ (.A1(_1020_),
    .A2(_1117_),
    .B(_1120_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3419_ (.A1(_1025_),
    .A2(_1118_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3420_ (.A1(_1024_),
    .A2(_1117_),
    .B(_1121_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3421_ (.A1(_1029_),
    .A2(_1118_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3422_ (.A1(_1028_),
    .A2(_1117_),
    .B(_1122_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3423_ (.I(_0961_),
    .Z(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3424_ (.A1(_0879_),
    .A2(_0933_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3425_ (.I(_1124_),
    .Z(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3426_ (.I(_1125_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3427_ (.I(_1124_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3428_ (.I(_1127_),
    .Z(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3429_ (.A1(_1037_),
    .A2(_1128_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3430_ (.A1(_1123_),
    .A2(_1126_),
    .B(_1129_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3431_ (.I(_0973_),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3432_ (.A1(_1041_),
    .A2(_1128_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3433_ (.A1(_1130_),
    .A2(_1126_),
    .B(_1131_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3434_ (.I(_0976_),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3435_ (.A1(_1043_),
    .A2(_1128_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3436_ (.A1(_1132_),
    .A2(_1126_),
    .B(_1133_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3437_ (.I(_0979_),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3438_ (.A1(_1045_),
    .A2(_1128_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3439_ (.A1(_1134_),
    .A2(_1126_),
    .B(_1135_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3440_ (.I(_1125_),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3441_ (.I(net28),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3442_ (.I(_1137_),
    .Z(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3443_ (.I(_1127_),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3444_ (.A1(_1138_),
    .A2(_1139_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3445_ (.A1(_1047_),
    .A2(_1136_),
    .B(_1140_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3446_ (.I(_0986_),
    .Z(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3447_ (.I(net29),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3448_ (.I(_1142_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3449_ (.A1(_1143_),
    .A2(_1139_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3450_ (.A1(_1141_),
    .A2(_1136_),
    .B(_1144_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3451_ (.I(_0990_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3452_ (.I(net30),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3453_ (.I(_1146_),
    .Z(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3454_ (.A1(_1147_),
    .A2(_1139_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3455_ (.A1(_1145_),
    .A2(_1136_),
    .B(_1148_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3456_ (.I(_0994_),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3457_ (.I(net31),
    .Z(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3458_ (.I(_1150_),
    .Z(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3459_ (.A1(_1151_),
    .A2(_1139_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3460_ (.A1(_1149_),
    .A2(_1136_),
    .B(_1152_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3461_ (.I(_0998_),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3462_ (.I(_1125_),
    .Z(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3463_ (.I(net32),
    .Z(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3464_ (.I(_1155_),
    .Z(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3465_ (.I(_1127_),
    .Z(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3466_ (.A1(_1156_),
    .A2(_1157_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3467_ (.A1(_1153_),
    .A2(_1154_),
    .B(_1158_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3468_ (.I(_1004_),
    .Z(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3469_ (.I(net33),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3470_ (.I(_1160_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3471_ (.A1(_1161_),
    .A2(_1157_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3472_ (.A1(_1159_),
    .A2(_1154_),
    .B(_1162_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3473_ (.I(_1008_),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3474_ (.A1(_1058_),
    .A2(_1157_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3475_ (.A1(_1163_),
    .A2(_1154_),
    .B(_1164_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3476_ (.I(net20),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3477_ (.I(_1165_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3478_ (.A1(_1166_),
    .A2(_1157_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3479_ (.A1(_1060_),
    .A2(_1154_),
    .B(_1167_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3480_ (.I(_1013_),
    .Z(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3481_ (.I(_1125_),
    .Z(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3482_ (.I(net21),
    .Z(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3483_ (.I(_1170_),
    .Z(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3484_ (.I(_1127_),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3485_ (.A1(_1171_),
    .A2(_1172_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3486_ (.A1(_1168_),
    .A2(_1169_),
    .B(_1173_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3487_ (.I(_1019_),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3488_ (.I(net22),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3489_ (.I(_1175_),
    .Z(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3490_ (.A1(_1176_),
    .A2(_1172_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3491_ (.A1(_1174_),
    .A2(_1169_),
    .B(_1177_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3492_ (.I(_1023_),
    .Z(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3493_ (.I(net23),
    .Z(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3494_ (.I(_1179_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3495_ (.A1(_1180_),
    .A2(_1172_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3496_ (.A1(_1178_),
    .A2(_1169_),
    .B(_1181_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3497_ (.I(_1027_),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3498_ (.I(net24),
    .Z(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3499_ (.I(_1183_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3500_ (.A1(_1184_),
    .A2(_1172_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3501_ (.A1(_1182_),
    .A2(_1169_),
    .B(_1185_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3502_ (.A1(_0930_),
    .A2(_0878_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3503_ (.A1(_1031_),
    .A2(_1186_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3504_ (.I(_1187_),
    .Z(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3505_ (.I(_1188_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3506_ (.I(net18),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3507_ (.I(_1190_),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3508_ (.I(_1187_),
    .Z(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3509_ (.I(_1192_),
    .Z(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3510_ (.A1(_1191_),
    .A2(_1193_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3511_ (.A1(_1123_),
    .A2(_1189_),
    .B(_1194_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3512_ (.I(net25),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3513_ (.I(_1195_),
    .Z(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3514_ (.A1(_1196_),
    .A2(_1193_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3515_ (.A1(_1130_),
    .A2(_1189_),
    .B(_1197_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3516_ (.I(net26),
    .Z(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3517_ (.I(_1198_),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3518_ (.A1(_1199_),
    .A2(_1193_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3519_ (.A1(_1132_),
    .A2(_1189_),
    .B(_1200_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3520_ (.I(net27),
    .Z(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3521_ (.I(_1201_),
    .Z(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3522_ (.A1(_1202_),
    .A2(_1193_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3523_ (.A1(_1134_),
    .A2(_1189_),
    .B(_1203_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3524_ (.I(_0794_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3525_ (.I(_1188_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3526_ (.I(_1192_),
    .Z(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3527_ (.A1(_1138_),
    .A2(_1206_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3528_ (.A1(_1204_),
    .A2(_1205_),
    .B(_1207_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3529_ (.A1(_1143_),
    .A2(_1206_),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3530_ (.A1(_1141_),
    .A2(_1205_),
    .B(_1208_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3531_ (.A1(_1147_),
    .A2(_1206_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3532_ (.A1(_1145_),
    .A2(_1205_),
    .B(_1209_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3533_ (.A1(_1151_),
    .A2(_1206_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3534_ (.A1(_1149_),
    .A2(_1205_),
    .B(_1210_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3535_ (.I(_1188_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3536_ (.I(_1192_),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3537_ (.A1(_1156_),
    .A2(_1212_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3538_ (.A1(_1153_),
    .A2(_1211_),
    .B(_1213_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3539_ (.A1(_1161_),
    .A2(_1212_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3540_ (.A1(_1159_),
    .A2(_1211_),
    .B(_1214_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3541_ (.I(net19),
    .Z(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3542_ (.I(_1215_),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3543_ (.A1(_1216_),
    .A2(_1212_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3544_ (.A1(_1163_),
    .A2(_1211_),
    .B(_1217_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3545_ (.I(_0821_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3546_ (.A1(_1166_),
    .A2(_1212_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3547_ (.A1(_1218_),
    .A2(_1211_),
    .B(_1219_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3548_ (.I(_1188_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3549_ (.I(_1192_),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3550_ (.A1(_1171_),
    .A2(_1221_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3551_ (.A1(_1168_),
    .A2(_1220_),
    .B(_1222_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3552_ (.A1(_1176_),
    .A2(_1221_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3553_ (.A1(_1174_),
    .A2(_1220_),
    .B(_1223_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3554_ (.A1(_1180_),
    .A2(_1221_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3555_ (.A1(_1178_),
    .A2(_1220_),
    .B(_1224_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3556_ (.A1(_1184_),
    .A2(_1221_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3557_ (.A1(_1182_),
    .A2(_1220_),
    .B(_1225_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3558_ (.A1(\Control_unit2.instr_stage2[8] ),
    .A2(_0751_),
    .A3(_0758_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3559_ (.A1(_0700_),
    .A2(_0764_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3560_ (.A1(_1227_),
    .A2(_0881_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3561_ (.I(_1228_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3562_ (.A1(_1226_),
    .A2(_1229_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3563_ (.I(_1230_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3564_ (.I(_1231_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3565_ (.I(_1230_),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3566_ (.I(_1233_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3567_ (.A1(_1191_),
    .A2(_1234_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3568_ (.A1(_1123_),
    .A2(_1232_),
    .B(_1235_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3569_ (.A1(_1196_),
    .A2(_1234_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3570_ (.A1(_1130_),
    .A2(_1232_),
    .B(_1236_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3571_ (.A1(_1199_),
    .A2(_1234_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3572_ (.A1(_1132_),
    .A2(_1232_),
    .B(_1237_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3573_ (.A1(_1202_),
    .A2(_1234_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3574_ (.A1(_1134_),
    .A2(_1232_),
    .B(_1238_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3575_ (.I(_1231_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3576_ (.I(_1233_),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3577_ (.A1(_1138_),
    .A2(_1240_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3578_ (.A1(_1204_),
    .A2(_1239_),
    .B(_1241_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3579_ (.A1(_1143_),
    .A2(_1240_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3580_ (.A1(_1141_),
    .A2(_1239_),
    .B(_1242_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3581_ (.A1(_1147_),
    .A2(_1240_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3582_ (.A1(_1145_),
    .A2(_1239_),
    .B(_1243_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3583_ (.A1(_1151_),
    .A2(_1240_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3584_ (.A1(_1149_),
    .A2(_1239_),
    .B(_1244_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3585_ (.I(_1231_),
    .Z(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3586_ (.I(_1233_),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3587_ (.A1(_1156_),
    .A2(_1246_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3588_ (.A1(_1153_),
    .A2(_1245_),
    .B(_1247_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3589_ (.A1(_1161_),
    .A2(_1246_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3590_ (.A1(_1159_),
    .A2(_1245_),
    .B(_1248_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3591_ (.A1(_1216_),
    .A2(_1246_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3592_ (.A1(_1163_),
    .A2(_1245_),
    .B(_1249_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3593_ (.A1(_1166_),
    .A2(_1246_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3594_ (.A1(_1218_),
    .A2(_1245_),
    .B(_1250_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3595_ (.I(_1231_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3596_ (.I(_1233_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3597_ (.A1(_1171_),
    .A2(_1252_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3598_ (.A1(_1168_),
    .A2(_1251_),
    .B(_1253_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3599_ (.A1(_1176_),
    .A2(_1252_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3600_ (.A1(_1174_),
    .A2(_1251_),
    .B(_1254_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3601_ (.A1(_1180_),
    .A2(_1252_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3602_ (.A1(_1178_),
    .A2(_1251_),
    .B(_1255_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3603_ (.A1(_1184_),
    .A2(_1252_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3604_ (.A1(_1182_),
    .A2(_1251_),
    .B(_1256_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3605_ (.A1(_0931_),
    .A2(_1229_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3606_ (.I(_1257_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3607_ (.I(_1258_),
    .Z(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3608_ (.I(_1257_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3609_ (.I(_1260_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3610_ (.A1(_1191_),
    .A2(_1261_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3611_ (.A1(_1123_),
    .A2(_1259_),
    .B(_1262_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3612_ (.A1(_1196_),
    .A2(_1261_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3613_ (.A1(_1130_),
    .A2(_1259_),
    .B(_1263_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3614_ (.A1(_1199_),
    .A2(_1261_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3615_ (.A1(_1132_),
    .A2(_1259_),
    .B(_1264_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3616_ (.A1(_1202_),
    .A2(_1261_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3617_ (.A1(_1134_),
    .A2(_1259_),
    .B(_1265_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3618_ (.I(_1258_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3619_ (.I(_1260_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3620_ (.A1(_1138_),
    .A2(_1267_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3621_ (.A1(_1204_),
    .A2(_1266_),
    .B(_1268_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3622_ (.A1(_1143_),
    .A2(_1267_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3623_ (.A1(_1141_),
    .A2(_1266_),
    .B(_1269_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3624_ (.A1(_1147_),
    .A2(_1267_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3625_ (.A1(_1145_),
    .A2(_1266_),
    .B(_1270_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3626_ (.A1(_1151_),
    .A2(_1267_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3627_ (.A1(_1149_),
    .A2(_1266_),
    .B(_1271_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3628_ (.I(_1258_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3629_ (.I(_1260_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3630_ (.A1(_1156_),
    .A2(_1273_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3631_ (.A1(_1153_),
    .A2(_1272_),
    .B(_1274_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3632_ (.A1(_1161_),
    .A2(_1273_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3633_ (.A1(_1159_),
    .A2(_1272_),
    .B(_1275_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3634_ (.A1(_1216_),
    .A2(_1273_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3635_ (.A1(_1163_),
    .A2(_1272_),
    .B(_1276_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3636_ (.A1(_1166_),
    .A2(_1273_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3637_ (.A1(_1218_),
    .A2(_1272_),
    .B(_1277_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3638_ (.I(_1258_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3639_ (.I(_1260_),
    .Z(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3640_ (.A1(_1171_),
    .A2(_1279_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3641_ (.A1(_1168_),
    .A2(_1278_),
    .B(_1280_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3642_ (.A1(_1176_),
    .A2(_1279_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3643_ (.A1(_1174_),
    .A2(_1278_),
    .B(_1281_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3644_ (.A1(_1180_),
    .A2(_1279_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3645_ (.A1(_1178_),
    .A2(_1278_),
    .B(_1282_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3646_ (.A1(_1184_),
    .A2(_1279_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3647_ (.A1(_1182_),
    .A2(_1278_),
    .B(_1283_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3648_ (.I(_2144_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3649_ (.I(_1284_),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3650_ (.A1(_0746_),
    .A2(_1032_),
    .A3(_0758_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3651_ (.A1(_1229_),
    .A2(_1286_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3652_ (.I(_1287_),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3653_ (.I(_1288_),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3654_ (.I(_1287_),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3655_ (.I(_1290_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3656_ (.A1(_1191_),
    .A2(_1291_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3657_ (.A1(_1285_),
    .A2(_1289_),
    .B(_1292_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3658_ (.I(_2170_),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3659_ (.I(_1293_),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3660_ (.A1(_1196_),
    .A2(_1291_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3661_ (.A1(_1294_),
    .A2(_1289_),
    .B(_1295_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3662_ (.I(_2188_),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3663_ (.I(_1296_),
    .Z(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3664_ (.A1(_1199_),
    .A2(_1291_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3665_ (.A1(_1297_),
    .A2(_1289_),
    .B(_1298_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3666_ (.I(_2210_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3667_ (.I(_1299_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3668_ (.A1(_1202_),
    .A2(_1291_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3669_ (.A1(_1300_),
    .A2(_1289_),
    .B(_1301_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3670_ (.I(_1288_),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3671_ (.I(_1137_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3672_ (.I(_1290_),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3673_ (.A1(_1303_),
    .A2(_1304_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3674_ (.A1(_1204_),
    .A2(_1302_),
    .B(_1305_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3675_ (.I(_2256_),
    .Z(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3676_ (.I(_1306_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3677_ (.I(_1142_),
    .Z(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3678_ (.A1(_1308_),
    .A2(_1304_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3679_ (.A1(_1307_),
    .A2(_1302_),
    .B(_1309_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3680_ (.I(_2277_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3681_ (.I(_1310_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3682_ (.I(_1146_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3683_ (.A1(_1312_),
    .A2(_1304_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3684_ (.A1(_1311_),
    .A2(_1302_),
    .B(_1313_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3685_ (.I(_2297_),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3686_ (.I(_1314_),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3687_ (.I(_1150_),
    .Z(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3688_ (.A1(_1316_),
    .A2(_1304_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3689_ (.A1(_1315_),
    .A2(_1302_),
    .B(_1317_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3690_ (.I(_2321_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3691_ (.I(_1318_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3692_ (.I(_1288_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3693_ (.I(_1155_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3694_ (.I(_1290_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3695_ (.A1(_1321_),
    .A2(_1322_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3696_ (.A1(_1319_),
    .A2(_1320_),
    .B(_1323_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3697_ (.I(_2334_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3698_ (.I(_1324_),
    .Z(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3699_ (.I(_1160_),
    .Z(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3700_ (.A1(_1326_),
    .A2(_1322_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3701_ (.A1(_1325_),
    .A2(_1320_),
    .B(_1327_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3702_ (.I(_2354_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3703_ (.I(_1328_),
    .Z(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3704_ (.A1(_1216_),
    .A2(_1322_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3705_ (.A1(_1329_),
    .A2(_1320_),
    .B(_1330_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3706_ (.I(_1165_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3707_ (.A1(_1331_),
    .A2(_1322_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3708_ (.A1(_1218_),
    .A2(_1320_),
    .B(_1332_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3709_ (.I(_0570_),
    .Z(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3710_ (.I(_1333_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3711_ (.I(_1288_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3712_ (.I(_1170_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3713_ (.I(_1290_),
    .Z(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3714_ (.A1(_1336_),
    .A2(_1337_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3715_ (.A1(_1334_),
    .A2(_1335_),
    .B(_1338_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3716_ (.I(_0591_),
    .Z(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3717_ (.I(_1339_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3718_ (.I(_1175_),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3719_ (.A1(_1341_),
    .A2(_1337_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3720_ (.A1(_1340_),
    .A2(_1335_),
    .B(_1342_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3721_ (.I(_0603_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3722_ (.I(_1343_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3723_ (.I(_1179_),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3724_ (.A1(_1345_),
    .A2(_1337_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3725_ (.A1(_1344_),
    .A2(_1335_),
    .B(_1346_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3726_ (.I(_0614_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3727_ (.I(_1347_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3728_ (.I(_1183_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3729_ (.A1(_1349_),
    .A2(_1337_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3730_ (.A1(_1348_),
    .A2(_1335_),
    .B(_1350_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3731_ (.A1(_1033_),
    .A2(_1229_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3732_ (.I(_1351_),
    .Z(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3733_ (.I(_1352_),
    .Z(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3734_ (.I(_1190_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3735_ (.I(_1351_),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3736_ (.I(_1355_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3737_ (.A1(_1354_),
    .A2(_1356_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3738_ (.A1(_1285_),
    .A2(_1353_),
    .B(_1357_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3739_ (.I(_1195_),
    .Z(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3740_ (.A1(_1358_),
    .A2(_1356_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3741_ (.A1(_1294_),
    .A2(_1353_),
    .B(_1359_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3742_ (.I(_1198_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3743_ (.A1(_1360_),
    .A2(_1356_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3744_ (.A1(_1297_),
    .A2(_1353_),
    .B(_1361_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3745_ (.I(_1201_),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3746_ (.A1(_1362_),
    .A2(_1356_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3747_ (.A1(_1300_),
    .A2(_1353_),
    .B(_1363_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3748_ (.I(_2232_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3749_ (.I(_1364_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3750_ (.I(_1352_),
    .Z(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3751_ (.I(_1355_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3752_ (.A1(_1303_),
    .A2(_1367_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3753_ (.A1(_1365_),
    .A2(_1366_),
    .B(_1368_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3754_ (.A1(_1308_),
    .A2(_1367_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3755_ (.A1(_1307_),
    .A2(_1366_),
    .B(_1369_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3756_ (.A1(_1312_),
    .A2(_1367_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3757_ (.A1(_1311_),
    .A2(_1366_),
    .B(_1370_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3758_ (.A1(_1316_),
    .A2(_1367_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3759_ (.A1(_1315_),
    .A2(_1366_),
    .B(_1371_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3760_ (.I(_1352_),
    .Z(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3761_ (.I(_1355_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3762_ (.A1(_1321_),
    .A2(_1373_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3763_ (.A1(_1319_),
    .A2(_1372_),
    .B(_1374_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3764_ (.A1(_1326_),
    .A2(_1373_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3765_ (.A1(_1325_),
    .A2(_1372_),
    .B(_1375_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3766_ (.I(_1215_),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3767_ (.A1(_1376_),
    .A2(_1373_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3768_ (.A1(_1329_),
    .A2(_1372_),
    .B(_1377_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3769_ (.I(_2370_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3770_ (.I(_1378_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3771_ (.A1(_1331_),
    .A2(_1373_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3772_ (.A1(_1379_),
    .A2(_1372_),
    .B(_1380_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3773_ (.I(_1352_),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3774_ (.I(_1355_),
    .Z(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3775_ (.A1(_1336_),
    .A2(_1382_),
    .ZN(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3776_ (.A1(_1334_),
    .A2(_1381_),
    .B(_1383_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3777_ (.A1(_1341_),
    .A2(_1382_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3778_ (.A1(_1340_),
    .A2(_1381_),
    .B(_1384_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3779_ (.A1(_1345_),
    .A2(_1382_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3780_ (.A1(_1344_),
    .A2(_1381_),
    .B(_1385_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3781_ (.A1(_1349_),
    .A2(_1382_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3782_ (.A1(_1348_),
    .A2(_1381_),
    .B(_1386_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3783_ (.A1(_0879_),
    .A2(_0966_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3784_ (.I(_1387_),
    .Z(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3785_ (.I(_1388_),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3786_ (.I(_1387_),
    .Z(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3787_ (.I(_1390_),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3788_ (.A1(_1354_),
    .A2(_1391_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3789_ (.A1(_1285_),
    .A2(_1389_),
    .B(_1392_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3790_ (.A1(_1358_),
    .A2(_1391_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3791_ (.A1(_1294_),
    .A2(_1389_),
    .B(_1393_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3792_ (.A1(_1360_),
    .A2(_1391_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3793_ (.A1(_1297_),
    .A2(_1389_),
    .B(_1394_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3794_ (.A1(_1362_),
    .A2(_1391_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3795_ (.A1(_1300_),
    .A2(_1389_),
    .B(_1395_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3796_ (.I(_1388_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3797_ (.I(_1390_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3798_ (.A1(_1303_),
    .A2(_1397_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3799_ (.A1(_1365_),
    .A2(_1396_),
    .B(_1398_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3800_ (.A1(_1308_),
    .A2(_1397_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3801_ (.A1(_1307_),
    .A2(_1396_),
    .B(_1399_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3802_ (.A1(_1312_),
    .A2(_1397_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3803_ (.A1(_1311_),
    .A2(_1396_),
    .B(_1400_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3804_ (.A1(_1316_),
    .A2(_1397_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3805_ (.A1(_1315_),
    .A2(_1396_),
    .B(_1401_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3806_ (.I(_1388_),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3807_ (.I(_1390_),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3808_ (.A1(_1321_),
    .A2(_1403_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3809_ (.A1(_1319_),
    .A2(_1402_),
    .B(_1404_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3810_ (.A1(_1326_),
    .A2(_1403_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3811_ (.A1(_1325_),
    .A2(_1402_),
    .B(_1405_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3812_ (.A1(_1376_),
    .A2(_1403_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3813_ (.A1(_1329_),
    .A2(_1402_),
    .B(_1406_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3814_ (.A1(_1331_),
    .A2(_1403_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3815_ (.A1(_1379_),
    .A2(_1402_),
    .B(_1407_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3816_ (.I(_1388_),
    .Z(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3817_ (.I(_1390_),
    .Z(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3818_ (.A1(_1336_),
    .A2(_1409_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3819_ (.A1(_1334_),
    .A2(_1408_),
    .B(_1410_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3820_ (.A1(_1341_),
    .A2(_1409_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3821_ (.A1(_1340_),
    .A2(_1408_),
    .B(_1411_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3822_ (.A1(_1345_),
    .A2(_1409_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3823_ (.A1(_1344_),
    .A2(_1408_),
    .B(_1412_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3824_ (.A1(_1349_),
    .A2(_1409_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3825_ (.A1(_1348_),
    .A2(_1408_),
    .B(_1413_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3826_ (.I(_1228_),
    .Z(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3827_ (.A1(_0964_),
    .A2(_1414_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3828_ (.I(_1415_),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3829_ (.I(_1416_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3830_ (.I(_1415_),
    .Z(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3831_ (.I(_1418_),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3832_ (.A1(_1354_),
    .A2(_1419_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3833_ (.A1(_1285_),
    .A2(_1417_),
    .B(_1420_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3834_ (.A1(_1358_),
    .A2(_1419_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3835_ (.A1(_1294_),
    .A2(_1417_),
    .B(_1421_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3836_ (.A1(_1360_),
    .A2(_1419_),
    .ZN(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3837_ (.A1(_1297_),
    .A2(_1417_),
    .B(_1422_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3838_ (.A1(_1362_),
    .A2(_1419_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3839_ (.A1(_1300_),
    .A2(_1417_),
    .B(_1423_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3840_ (.I(_1416_),
    .Z(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3841_ (.I(_1418_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3842_ (.A1(_1303_),
    .A2(_1425_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3843_ (.A1(_1365_),
    .A2(_1424_),
    .B(_1426_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3844_ (.A1(_1308_),
    .A2(_1425_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3845_ (.A1(_1307_),
    .A2(_1424_),
    .B(_1427_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3846_ (.A1(_1312_),
    .A2(_1425_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3847_ (.A1(_1311_),
    .A2(_1424_),
    .B(_1428_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3848_ (.A1(_1316_),
    .A2(_1425_),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3849_ (.A1(_1315_),
    .A2(_1424_),
    .B(_1429_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3850_ (.I(_1416_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3851_ (.I(_1418_),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3852_ (.A1(_1321_),
    .A2(_1431_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3853_ (.A1(_1319_),
    .A2(_1430_),
    .B(_1432_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3854_ (.A1(_1326_),
    .A2(_1431_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3855_ (.A1(_1325_),
    .A2(_1430_),
    .B(_1433_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3856_ (.A1(_1376_),
    .A2(_1431_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3857_ (.A1(_1329_),
    .A2(_1430_),
    .B(_1434_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3858_ (.A1(_1331_),
    .A2(_1431_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3859_ (.A1(_1379_),
    .A2(_1430_),
    .B(_1435_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3860_ (.I(_1416_),
    .Z(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3861_ (.I(_1418_),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3862_ (.A1(_1336_),
    .A2(_1437_),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3863_ (.A1(_1334_),
    .A2(_1436_),
    .B(_1438_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3864_ (.A1(_1341_),
    .A2(_1437_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3865_ (.A1(_1340_),
    .A2(_1436_),
    .B(_1439_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3866_ (.A1(_1345_),
    .A2(_1437_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3867_ (.A1(_1344_),
    .A2(_1436_),
    .B(_1440_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3868_ (.A1(_1349_),
    .A2(_1437_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3869_ (.A1(_1348_),
    .A2(_1436_),
    .B(_1441_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3870_ (.I(_1284_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3871_ (.A1(_0879_),
    .A2(_1414_),
    .ZN(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3872_ (.I(_1443_),
    .Z(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3873_ (.I(_1444_),
    .Z(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3874_ (.I(_1443_),
    .Z(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3875_ (.I(_1446_),
    .Z(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3876_ (.A1(_1354_),
    .A2(_1447_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3877_ (.A1(_1442_),
    .A2(_1445_),
    .B(_1448_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3878_ (.I(_1293_),
    .Z(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3879_ (.A1(_1358_),
    .A2(_1447_),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3880_ (.A1(_1449_),
    .A2(_1445_),
    .B(_1450_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3881_ (.I(_1296_),
    .Z(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3882_ (.A1(_1360_),
    .A2(_1447_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3883_ (.A1(_1451_),
    .A2(_1445_),
    .B(_1452_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3884_ (.I(_1299_),
    .Z(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3885_ (.A1(_1362_),
    .A2(_1447_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3886_ (.A1(_1453_),
    .A2(_1445_),
    .B(_1454_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3887_ (.I(_1444_),
    .Z(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3888_ (.I(_1137_),
    .Z(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3889_ (.I(_1446_),
    .Z(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3890_ (.A1(_1456_),
    .A2(_1457_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3891_ (.A1(_1365_),
    .A2(_1455_),
    .B(_1458_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3892_ (.I(_1306_),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3893_ (.I(_1142_),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3894_ (.A1(_1460_),
    .A2(_1457_),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3895_ (.A1(_1459_),
    .A2(_1455_),
    .B(_1461_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3896_ (.I(_1310_),
    .Z(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3897_ (.I(_1146_),
    .Z(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3898_ (.A1(_1463_),
    .A2(_1457_),
    .ZN(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3899_ (.A1(_1462_),
    .A2(_1455_),
    .B(_1464_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3900_ (.I(_1314_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3901_ (.I(_1150_),
    .Z(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3902_ (.A1(_1466_),
    .A2(_1457_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3903_ (.A1(_1465_),
    .A2(_1455_),
    .B(_1467_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3904_ (.I(_1318_),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3905_ (.I(_1444_),
    .Z(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3906_ (.I(_1155_),
    .Z(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3907_ (.I(_1446_),
    .Z(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3908_ (.A1(_1470_),
    .A2(_1471_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3909_ (.A1(_1468_),
    .A2(_1469_),
    .B(_1472_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3910_ (.I(_1324_),
    .Z(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3911_ (.I(_1160_),
    .Z(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3912_ (.A1(_1474_),
    .A2(_1471_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3913_ (.A1(_1473_),
    .A2(_1469_),
    .B(_1475_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3914_ (.I(_1328_),
    .Z(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3915_ (.A1(_1376_),
    .A2(_1471_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3916_ (.A1(_1476_),
    .A2(_1469_),
    .B(_1477_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3917_ (.I(_1165_),
    .Z(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3918_ (.A1(_1478_),
    .A2(_1471_),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3919_ (.A1(_1379_),
    .A2(_1469_),
    .B(_1479_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3920_ (.I(_1333_),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3921_ (.I(_1444_),
    .Z(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3922_ (.I(_1170_),
    .Z(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3923_ (.I(_1446_),
    .Z(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3924_ (.A1(_1482_),
    .A2(_1483_),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3925_ (.A1(_1480_),
    .A2(_1481_),
    .B(_1484_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3926_ (.I(_1339_),
    .Z(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3927_ (.I(_1175_),
    .Z(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3928_ (.A1(_1486_),
    .A2(_1483_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3929_ (.A1(_1485_),
    .A2(_1481_),
    .B(_1487_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3930_ (.I(_1343_),
    .Z(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3931_ (.I(_1179_),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3932_ (.A1(_1489_),
    .A2(_1483_),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3933_ (.A1(_1488_),
    .A2(_1481_),
    .B(_1490_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3934_ (.I(_1347_),
    .Z(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3935_ (.I(_1183_),
    .Z(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3936_ (.A1(_1492_),
    .A2(_1483_),
    .ZN(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3937_ (.A1(_1491_),
    .A2(_1481_),
    .B(_1493_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3938_ (.A1(_1186_),
    .A2(_1414_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3939_ (.I(_1494_),
    .Z(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3940_ (.I(_1495_),
    .Z(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3941_ (.I(_1190_),
    .Z(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3942_ (.I(_1494_),
    .Z(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3943_ (.I(_1498_),
    .Z(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3944_ (.A1(_1497_),
    .A2(_1499_),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3945_ (.A1(_1442_),
    .A2(_1496_),
    .B(_1500_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3946_ (.I(_1195_),
    .Z(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3947_ (.A1(_1501_),
    .A2(_1499_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3948_ (.A1(_1449_),
    .A2(_1496_),
    .B(_1502_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3949_ (.I(_1198_),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3950_ (.A1(_1503_),
    .A2(_1499_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3951_ (.A1(_1451_),
    .A2(_1496_),
    .B(_1504_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3952_ (.I(_1201_),
    .Z(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3953_ (.A1(_1505_),
    .A2(_1499_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3954_ (.A1(_1453_),
    .A2(_1496_),
    .B(_1506_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3955_ (.I(_1364_),
    .Z(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3956_ (.I(_1495_),
    .Z(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3957_ (.I(_1498_),
    .Z(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3958_ (.A1(_1456_),
    .A2(_1509_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3959_ (.A1(_1507_),
    .A2(_1508_),
    .B(_1510_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3960_ (.A1(_1460_),
    .A2(_1509_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3961_ (.A1(_1459_),
    .A2(_1508_),
    .B(_1511_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3962_ (.A1(_1463_),
    .A2(_1509_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3963_ (.A1(_1462_),
    .A2(_1508_),
    .B(_1512_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3964_ (.A1(_1466_),
    .A2(_1509_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3965_ (.A1(_1465_),
    .A2(_1508_),
    .B(_1513_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3966_ (.I(_1495_),
    .Z(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3967_ (.I(_1498_),
    .Z(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3968_ (.A1(_1470_),
    .A2(_1515_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3969_ (.A1(_1468_),
    .A2(_1514_),
    .B(_1516_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3970_ (.A1(_1474_),
    .A2(_1515_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3971_ (.A1(_1473_),
    .A2(_1514_),
    .B(_1517_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3972_ (.I(_1215_),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3973_ (.A1(_1518_),
    .A2(_1515_),
    .ZN(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3974_ (.A1(_1476_),
    .A2(_1514_),
    .B(_1519_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3975_ (.I(_1378_),
    .Z(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3976_ (.A1(_1478_),
    .A2(_1515_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3977_ (.A1(_1520_),
    .A2(_1514_),
    .B(_1521_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3978_ (.I(_1495_),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3979_ (.I(_1498_),
    .Z(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3980_ (.A1(_1482_),
    .A2(_1523_),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3981_ (.A1(_1480_),
    .A2(_1522_),
    .B(_1524_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3982_ (.A1(_1486_),
    .A2(_1523_),
    .ZN(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3983_ (.A1(_1485_),
    .A2(_1522_),
    .B(_1525_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3984_ (.A1(_1489_),
    .A2(_1523_),
    .ZN(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3985_ (.A1(_1488_),
    .A2(_1522_),
    .B(_1526_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3986_ (.A1(_1492_),
    .A2(_1523_),
    .ZN(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3987_ (.A1(_1491_),
    .A2(_1522_),
    .B(_1527_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3988_ (.I(_0882_),
    .Z(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3989_ (.A1(_1528_),
    .A2(_1226_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3990_ (.I(_1529_),
    .Z(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3991_ (.I(_1530_),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3992_ (.I(_1529_),
    .Z(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3993_ (.I(_1532_),
    .Z(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3994_ (.A1(_1497_),
    .A2(_1533_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3995_ (.A1(_1442_),
    .A2(_1531_),
    .B(_1534_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3996_ (.A1(_1501_),
    .A2(_1533_),
    .ZN(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3997_ (.A1(_1449_),
    .A2(_1531_),
    .B(_1535_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3998_ (.A1(_1503_),
    .A2(_1533_),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3999_ (.A1(_1451_),
    .A2(_1531_),
    .B(_1536_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4000_ (.A1(_1505_),
    .A2(_1533_),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4001_ (.A1(_1453_),
    .A2(_1531_),
    .B(_1537_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4002_ (.I(_1530_),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4003_ (.I(_1532_),
    .Z(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4004_ (.A1(_1456_),
    .A2(_1539_),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4005_ (.A1(_1507_),
    .A2(_1538_),
    .B(_1540_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4006_ (.A1(_1460_),
    .A2(_1539_),
    .ZN(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4007_ (.A1(_1459_),
    .A2(_1538_),
    .B(_1541_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4008_ (.A1(_1463_),
    .A2(_1539_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4009_ (.A1(_1462_),
    .A2(_1538_),
    .B(_1542_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4010_ (.A1(_1466_),
    .A2(_1539_),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4011_ (.A1(_1465_),
    .A2(_1538_),
    .B(_1543_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4012_ (.I(_1530_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4013_ (.I(_1532_),
    .Z(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4014_ (.A1(_1470_),
    .A2(_1545_),
    .ZN(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4015_ (.A1(_1468_),
    .A2(_1544_),
    .B(_1546_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4016_ (.A1(_1474_),
    .A2(_1545_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4017_ (.A1(_1473_),
    .A2(_1544_),
    .B(_1547_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4018_ (.A1(_1518_),
    .A2(_1545_),
    .ZN(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4019_ (.A1(_1476_),
    .A2(_1544_),
    .B(_1548_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4020_ (.A1(_1478_),
    .A2(_1545_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4021_ (.A1(_1520_),
    .A2(_1544_),
    .B(_1549_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4022_ (.I(_1530_),
    .Z(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4023_ (.I(_1532_),
    .Z(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4024_ (.A1(_1482_),
    .A2(_1551_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4025_ (.A1(_1480_),
    .A2(_1550_),
    .B(_1552_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4026_ (.A1(_1486_),
    .A2(_1551_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4027_ (.A1(_1485_),
    .A2(_1550_),
    .B(_1553_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4028_ (.A1(_1489_),
    .A2(_1551_),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4029_ (.A1(_1488_),
    .A2(_1550_),
    .B(_1554_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4030_ (.A1(_1492_),
    .A2(_1551_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4031_ (.A1(_1491_),
    .A2(_1550_),
    .B(_1555_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4032_ (.A1(_1528_),
    .A2(_0931_),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4033_ (.I(_1556_),
    .Z(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4034_ (.I(_1557_),
    .Z(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4035_ (.I(_1556_),
    .Z(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4036_ (.I(_1559_),
    .Z(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4037_ (.A1(_1497_),
    .A2(_1560_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4038_ (.A1(_1442_),
    .A2(_1558_),
    .B(_1561_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4039_ (.A1(_1501_),
    .A2(_1560_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4040_ (.A1(_1449_),
    .A2(_1558_),
    .B(_1562_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4041_ (.A1(_1503_),
    .A2(_1560_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4042_ (.A1(_1451_),
    .A2(_1558_),
    .B(_1563_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4043_ (.A1(_1505_),
    .A2(_1560_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4044_ (.A1(_1453_),
    .A2(_1558_),
    .B(_1564_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4045_ (.I(_1557_),
    .Z(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4046_ (.I(_1559_),
    .Z(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4047_ (.A1(_1456_),
    .A2(_1566_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4048_ (.A1(_1507_),
    .A2(_1565_),
    .B(_1567_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4049_ (.A1(_1460_),
    .A2(_1566_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4050_ (.A1(_1459_),
    .A2(_1565_),
    .B(_1568_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4051_ (.A1(_1463_),
    .A2(_1566_),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4052_ (.A1(_1462_),
    .A2(_1565_),
    .B(_1569_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4053_ (.A1(_1466_),
    .A2(_1566_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4054_ (.A1(_1465_),
    .A2(_1565_),
    .B(_1570_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4055_ (.I(_1557_),
    .Z(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4056_ (.I(_1559_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4057_ (.A1(_1470_),
    .A2(_1572_),
    .ZN(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4058_ (.A1(_1468_),
    .A2(_1571_),
    .B(_1573_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4059_ (.A1(_1474_),
    .A2(_1572_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4060_ (.A1(_1473_),
    .A2(_1571_),
    .B(_1574_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4061_ (.A1(_1518_),
    .A2(_1572_),
    .ZN(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4062_ (.A1(_1476_),
    .A2(_1571_),
    .B(_1575_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4063_ (.A1(_1478_),
    .A2(_1572_),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4064_ (.A1(_1520_),
    .A2(_1571_),
    .B(_1576_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4065_ (.I(_1557_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4066_ (.I(_1559_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4067_ (.A1(_1482_),
    .A2(_1578_),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4068_ (.A1(_1480_),
    .A2(_1577_),
    .B(_1579_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4069_ (.A1(_1486_),
    .A2(_1578_),
    .ZN(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4070_ (.A1(_1485_),
    .A2(_1577_),
    .B(_1580_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4071_ (.A1(_1489_),
    .A2(_1578_),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4072_ (.A1(_1488_),
    .A2(_1577_),
    .B(_1581_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4073_ (.A1(_1492_),
    .A2(_1578_),
    .ZN(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4074_ (.A1(_1491_),
    .A2(_1577_),
    .B(_1582_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4075_ (.I(_1284_),
    .Z(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4076_ (.A1(_1528_),
    .A2(_1286_),
    .ZN(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4077_ (.I(_1584_),
    .Z(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4078_ (.I(_1585_),
    .Z(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4079_ (.I(_1584_),
    .Z(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4080_ (.I(_1587_),
    .Z(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4081_ (.A1(_1497_),
    .A2(_1588_),
    .ZN(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4082_ (.A1(_1583_),
    .A2(_1586_),
    .B(_1589_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4083_ (.I(_1293_),
    .Z(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4084_ (.A1(_1501_),
    .A2(_1588_),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4085_ (.A1(_1590_),
    .A2(_1586_),
    .B(_1591_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4086_ (.I(_1296_),
    .Z(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4087_ (.A1(_1503_),
    .A2(_1588_),
    .ZN(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4088_ (.A1(_1592_),
    .A2(_1586_),
    .B(_1593_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4089_ (.I(_1299_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4090_ (.A1(_1505_),
    .A2(_1588_),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4091_ (.A1(_1594_),
    .A2(_1586_),
    .B(_1595_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4092_ (.I(_1585_),
    .Z(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4093_ (.I(_1137_),
    .Z(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4094_ (.I(_1587_),
    .Z(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4095_ (.A1(_1597_),
    .A2(_1598_),
    .ZN(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4096_ (.A1(_1507_),
    .A2(_1596_),
    .B(_1599_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4097_ (.I(_1306_),
    .Z(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4098_ (.I(_1142_),
    .Z(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4099_ (.A1(_1601_),
    .A2(_1598_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4100_ (.A1(_1600_),
    .A2(_1596_),
    .B(_1602_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4101_ (.I(_1310_),
    .Z(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4102_ (.I(_1146_),
    .Z(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4103_ (.A1(_1604_),
    .A2(_1598_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4104_ (.A1(_1603_),
    .A2(_1596_),
    .B(_1605_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4105_ (.I(_1314_),
    .Z(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4106_ (.I(_1150_),
    .Z(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4107_ (.A1(_1607_),
    .A2(_1598_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4108_ (.A1(_1606_),
    .A2(_1596_),
    .B(_1608_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4109_ (.I(_1318_),
    .Z(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4110_ (.I(_1585_),
    .Z(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4111_ (.I(_1155_),
    .Z(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4112_ (.I(_1587_),
    .Z(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4113_ (.A1(_1611_),
    .A2(_1612_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4114_ (.A1(_1609_),
    .A2(_1610_),
    .B(_1613_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4115_ (.I(_1324_),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4116_ (.I(_1160_),
    .Z(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4117_ (.A1(_1615_),
    .A2(_1612_),
    .ZN(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4118_ (.A1(_1614_),
    .A2(_1610_),
    .B(_1616_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4119_ (.I(_1328_),
    .Z(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4120_ (.A1(_1518_),
    .A2(_1612_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4121_ (.A1(_1617_),
    .A2(_1610_),
    .B(_1618_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4122_ (.I(_1165_),
    .Z(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4123_ (.A1(_1619_),
    .A2(_1612_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4124_ (.A1(_1520_),
    .A2(_1610_),
    .B(_1620_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4125_ (.I(_1333_),
    .Z(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4126_ (.I(_1585_),
    .Z(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4127_ (.I(_1170_),
    .Z(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4128_ (.I(_1587_),
    .Z(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4129_ (.A1(_1623_),
    .A2(_1624_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4130_ (.A1(_1621_),
    .A2(_1622_),
    .B(_1625_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4131_ (.I(_1339_),
    .Z(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4132_ (.I(_1175_),
    .Z(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4133_ (.A1(_1627_),
    .A2(_1624_),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4134_ (.A1(_1626_),
    .A2(_1622_),
    .B(_1628_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4135_ (.I(_1343_),
    .Z(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4136_ (.I(_1179_),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4137_ (.A1(_1630_),
    .A2(_1624_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4138_ (.A1(_1629_),
    .A2(_1622_),
    .B(_1631_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4139_ (.I(_1347_),
    .Z(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4140_ (.I(_1183_),
    .Z(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4141_ (.A1(_1633_),
    .A2(_1624_),
    .ZN(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4142_ (.A1(_1632_),
    .A2(_1622_),
    .B(_1634_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4143_ (.A1(_1528_),
    .A2(_1033_),
    .ZN(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4144_ (.I(_1635_),
    .Z(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4145_ (.I(_1636_),
    .Z(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4146_ (.I(_1190_),
    .Z(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4147_ (.I(_1635_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4148_ (.I(_1639_),
    .Z(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4149_ (.A1(_1638_),
    .A2(_1640_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4150_ (.A1(_1583_),
    .A2(_1637_),
    .B(_1641_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4151_ (.I(_1195_),
    .Z(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4152_ (.A1(_1642_),
    .A2(_1640_),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4153_ (.A1(_1590_),
    .A2(_1637_),
    .B(_1643_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4154_ (.I(_1198_),
    .Z(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4155_ (.A1(_1644_),
    .A2(_1640_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4156_ (.A1(_1592_),
    .A2(_1637_),
    .B(_1645_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4157_ (.I(_1201_),
    .Z(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4158_ (.A1(_1646_),
    .A2(_1640_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4159_ (.A1(_1594_),
    .A2(_1637_),
    .B(_1647_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4160_ (.I(_1364_),
    .Z(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4161_ (.I(_1636_),
    .Z(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4162_ (.I(_1639_),
    .Z(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4163_ (.A1(_1597_),
    .A2(_1650_),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4164_ (.A1(_1648_),
    .A2(_1649_),
    .B(_1651_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4165_ (.A1(_1601_),
    .A2(_1650_),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4166_ (.A1(_1600_),
    .A2(_1649_),
    .B(_1652_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4167_ (.A1(_1604_),
    .A2(_1650_),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4168_ (.A1(_1603_),
    .A2(_1649_),
    .B(_1653_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4169_ (.A1(_1607_),
    .A2(_1650_),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4170_ (.A1(_1606_),
    .A2(_1649_),
    .B(_1654_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4171_ (.I(_1636_),
    .Z(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4172_ (.I(_1639_),
    .Z(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4173_ (.A1(_1611_),
    .A2(_1656_),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4174_ (.A1(_1609_),
    .A2(_1655_),
    .B(_1657_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4175_ (.A1(_1615_),
    .A2(_1656_),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4176_ (.A1(_1614_),
    .A2(_1655_),
    .B(_1658_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4177_ (.I(_1215_),
    .Z(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4178_ (.A1(_1659_),
    .A2(_1656_),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4179_ (.A1(_1617_),
    .A2(_1655_),
    .B(_1660_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4180_ (.I(_1378_),
    .Z(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4181_ (.A1(_1619_),
    .A2(_1656_),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4182_ (.A1(_1661_),
    .A2(_1655_),
    .B(_1662_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4183_ (.I(_1636_),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4184_ (.I(_1639_),
    .Z(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4185_ (.A1(_1623_),
    .A2(_1664_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4186_ (.A1(_1621_),
    .A2(_1663_),
    .B(_1665_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4187_ (.A1(_1627_),
    .A2(_1664_),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4188_ (.A1(_1626_),
    .A2(_1663_),
    .B(_1666_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4189_ (.A1(_1630_),
    .A2(_1664_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4190_ (.A1(_1629_),
    .A2(_1663_),
    .B(_1667_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4191_ (.A1(_1633_),
    .A2(_1664_),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4192_ (.A1(_1632_),
    .A2(_1663_),
    .B(_1668_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4193_ (.A1(_0883_),
    .A2(_1068_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4194_ (.I(_1669_),
    .Z(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4195_ (.I(_1670_),
    .Z(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4196_ (.I(_1669_),
    .Z(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4197_ (.I(_1672_),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4198_ (.A1(_1638_),
    .A2(_1673_),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4199_ (.A1(_1583_),
    .A2(_1671_),
    .B(_1674_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4200_ (.A1(_1642_),
    .A2(_1673_),
    .ZN(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4201_ (.A1(_1590_),
    .A2(_1671_),
    .B(_1675_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4202_ (.A1(_1644_),
    .A2(_1673_),
    .ZN(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4203_ (.A1(_1592_),
    .A2(_1671_),
    .B(_1676_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4204_ (.A1(_1646_),
    .A2(_1673_),
    .ZN(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4205_ (.A1(_1594_),
    .A2(_1671_),
    .B(_1677_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4206_ (.I(_1670_),
    .Z(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4207_ (.I(_1672_),
    .Z(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4208_ (.A1(_1597_),
    .A2(_1679_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4209_ (.A1(_1648_),
    .A2(_1678_),
    .B(_1680_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4210_ (.A1(_1601_),
    .A2(_1679_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4211_ (.A1(_1600_),
    .A2(_1678_),
    .B(_1681_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4212_ (.A1(_1604_),
    .A2(_1679_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4213_ (.A1(_1603_),
    .A2(_1678_),
    .B(_1682_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4214_ (.A1(_1607_),
    .A2(_1679_),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4215_ (.A1(_1606_),
    .A2(_1678_),
    .B(_1683_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4216_ (.I(_1670_),
    .Z(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4217_ (.I(_1672_),
    .Z(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4218_ (.A1(_1611_),
    .A2(_1685_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4219_ (.A1(_1609_),
    .A2(_1684_),
    .B(_1686_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4220_ (.A1(_1615_),
    .A2(_1685_),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4221_ (.A1(_1614_),
    .A2(_1684_),
    .B(_1687_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4222_ (.A1(_1659_),
    .A2(_1685_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4223_ (.A1(_1617_),
    .A2(_1684_),
    .B(_1688_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4224_ (.A1(_1619_),
    .A2(_1685_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4225_ (.A1(_1661_),
    .A2(_1684_),
    .B(_1689_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4226_ (.I(_1670_),
    .Z(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4227_ (.I(_1672_),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4228_ (.A1(_1623_),
    .A2(_1691_),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4229_ (.A1(_1621_),
    .A2(_1690_),
    .B(_1692_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4230_ (.A1(_1627_),
    .A2(_1691_),
    .ZN(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4231_ (.A1(_1626_),
    .A2(_1690_),
    .B(_1693_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4232_ (.A1(_1630_),
    .A2(_1691_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4233_ (.A1(_1629_),
    .A2(_1690_),
    .B(_1694_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4234_ (.A1(_1633_),
    .A2(_1691_),
    .ZN(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4235_ (.A1(_1632_),
    .A2(_1690_),
    .B(_1695_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4236_ (.A1(_0883_),
    .A2(_0964_),
    .ZN(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4237_ (.I(_1696_),
    .Z(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4238_ (.I(_1697_),
    .Z(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4239_ (.I(_1696_),
    .Z(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4240_ (.I(_1699_),
    .Z(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4241_ (.A1(_1638_),
    .A2(_1700_),
    .ZN(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4242_ (.A1(_1583_),
    .A2(_1698_),
    .B(_1701_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4243_ (.A1(_1642_),
    .A2(_1700_),
    .ZN(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4244_ (.A1(_1590_),
    .A2(_1698_),
    .B(_1702_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4245_ (.A1(_1644_),
    .A2(_1700_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4246_ (.A1(_1592_),
    .A2(_1698_),
    .B(_1703_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4247_ (.A1(_1646_),
    .A2(_1700_),
    .ZN(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4248_ (.A1(_1594_),
    .A2(_1698_),
    .B(_1704_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4249_ (.I(_1697_),
    .Z(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4250_ (.I(_1699_),
    .Z(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4251_ (.A1(_1597_),
    .A2(_1706_),
    .ZN(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4252_ (.A1(_1648_),
    .A2(_1705_),
    .B(_1707_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4253_ (.A1(_1601_),
    .A2(_1706_),
    .ZN(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4254_ (.A1(_1600_),
    .A2(_1705_),
    .B(_1708_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4255_ (.A1(_1604_),
    .A2(_1706_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4256_ (.A1(_1603_),
    .A2(_1705_),
    .B(_1709_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4257_ (.A1(_1607_),
    .A2(_1706_),
    .ZN(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4258_ (.A1(_1606_),
    .A2(_1705_),
    .B(_1710_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4259_ (.I(_1697_),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4260_ (.I(_1699_),
    .Z(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4261_ (.A1(_1611_),
    .A2(_1712_),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4262_ (.A1(_1609_),
    .A2(_1711_),
    .B(_1713_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4263_ (.A1(_1615_),
    .A2(_1712_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4264_ (.A1(_1614_),
    .A2(_1711_),
    .B(_1714_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4265_ (.A1(_1659_),
    .A2(_1712_),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4266_ (.A1(_1617_),
    .A2(_1711_),
    .B(_1715_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4267_ (.A1(_1619_),
    .A2(_1712_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4268_ (.A1(_1661_),
    .A2(_1711_),
    .B(_1716_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4269_ (.I(_1697_),
    .Z(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4270_ (.I(_1699_),
    .Z(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4271_ (.A1(_1623_),
    .A2(_1718_),
    .ZN(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4272_ (.A1(_1621_),
    .A2(_1717_),
    .B(_1719_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4273_ (.A1(_1627_),
    .A2(_1718_),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4274_ (.A1(_1626_),
    .A2(_1717_),
    .B(_1720_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4275_ (.A1(_1630_),
    .A2(_1718_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4276_ (.A1(_1629_),
    .A2(_1717_),
    .B(_1721_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4277_ (.A1(_1633_),
    .A2(_1718_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4278_ (.A1(_1632_),
    .A2(_1717_),
    .B(_1722_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4279_ (.I(_1284_),
    .Z(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4280_ (.I(_0965_),
    .Z(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4281_ (.A1(_1724_),
    .A2(_1186_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4282_ (.I(_1725_),
    .Z(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4283_ (.I(_1726_),
    .Z(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4284_ (.I(_1725_),
    .Z(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4285_ (.I(_1728_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4286_ (.A1(_1638_),
    .A2(_1729_),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4287_ (.A1(_1723_),
    .A2(_1727_),
    .B(_1730_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4288_ (.I(_1293_),
    .Z(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4289_ (.A1(_1642_),
    .A2(_1729_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4290_ (.A1(_1731_),
    .A2(_1727_),
    .B(_1732_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4291_ (.I(_1296_),
    .Z(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4292_ (.A1(_1644_),
    .A2(_1729_),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4293_ (.A1(_1733_),
    .A2(_1727_),
    .B(_1734_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4294_ (.I(_1299_),
    .Z(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4295_ (.A1(_1646_),
    .A2(_1729_),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4296_ (.A1(_1735_),
    .A2(_1727_),
    .B(_1736_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4297_ (.I(_1726_),
    .Z(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4298_ (.I(net28),
    .Z(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4299_ (.I(_1728_),
    .Z(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4300_ (.A1(_1738_),
    .A2(_1739_),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4301_ (.A1(_1648_),
    .A2(_1737_),
    .B(_1740_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4302_ (.I(_1306_),
    .Z(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4303_ (.I(net29),
    .Z(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4304_ (.A1(_1742_),
    .A2(_1739_),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4305_ (.A1(_1741_),
    .A2(_1737_),
    .B(_1743_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4306_ (.I(_1310_),
    .Z(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4307_ (.I(net30),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4308_ (.A1(_1745_),
    .A2(_1739_),
    .ZN(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4309_ (.A1(_1744_),
    .A2(_1737_),
    .B(_1746_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4310_ (.I(_1314_),
    .Z(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4311_ (.I(net31),
    .Z(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4312_ (.A1(_1748_),
    .A2(_1739_),
    .ZN(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4313_ (.A1(_1747_),
    .A2(_1737_),
    .B(_1749_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4314_ (.I(_1318_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4315_ (.I(_1726_),
    .Z(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4316_ (.I(net32),
    .Z(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4317_ (.I(_1728_),
    .Z(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4318_ (.A1(_1752_),
    .A2(_1753_),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4319_ (.A1(_1750_),
    .A2(_1751_),
    .B(_1754_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4320_ (.I(_1324_),
    .Z(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4321_ (.I(net33),
    .Z(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4322_ (.A1(_1756_),
    .A2(_1753_),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4323_ (.A1(_1755_),
    .A2(_1751_),
    .B(_1757_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4324_ (.I(_1328_),
    .Z(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4325_ (.A1(_1659_),
    .A2(_1753_),
    .ZN(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4326_ (.A1(_1758_),
    .A2(_1751_),
    .B(_1759_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4327_ (.I(net20),
    .Z(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4328_ (.A1(_1760_),
    .A2(_1753_),
    .ZN(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4329_ (.A1(_1661_),
    .A2(_1751_),
    .B(_1761_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4330_ (.I(_1333_),
    .Z(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4331_ (.I(_1726_),
    .Z(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4332_ (.I(net21),
    .Z(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4333_ (.I(_1728_),
    .Z(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4334_ (.A1(_1764_),
    .A2(_1765_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4335_ (.A1(_1762_),
    .A2(_1763_),
    .B(_1766_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4336_ (.I(_1339_),
    .Z(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4337_ (.I(net22),
    .Z(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4338_ (.A1(_1768_),
    .A2(_1765_),
    .ZN(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4339_ (.A1(_1767_),
    .A2(_1763_),
    .B(_1769_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4340_ (.I(_1343_),
    .Z(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4341_ (.I(net23),
    .Z(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4342_ (.A1(_1771_),
    .A2(_1765_),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4343_ (.A1(_1770_),
    .A2(_1763_),
    .B(_1772_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4344_ (.I(_1347_),
    .Z(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4345_ (.I(net24),
    .Z(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4346_ (.A1(_1774_),
    .A2(_1765_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4347_ (.A1(_1773_),
    .A2(_1763_),
    .B(_1775_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4348_ (.A1(_0883_),
    .A2(_1186_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4349_ (.I(_1776_),
    .Z(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4350_ (.I(_1777_),
    .Z(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4351_ (.I(net18),
    .Z(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4352_ (.I(_1776_),
    .Z(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4353_ (.I(_1780_),
    .Z(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4354_ (.A1(_1779_),
    .A2(_1781_),
    .ZN(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4355_ (.A1(_1723_),
    .A2(_1778_),
    .B(_1782_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4356_ (.I(net25),
    .Z(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4357_ (.A1(_1783_),
    .A2(_1781_),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4358_ (.A1(_1731_),
    .A2(_1778_),
    .B(_1784_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4359_ (.I(net26),
    .Z(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4360_ (.A1(_1785_),
    .A2(_1781_),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4361_ (.A1(_1733_),
    .A2(_1778_),
    .B(_1786_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4362_ (.I(net27),
    .Z(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4363_ (.A1(_1787_),
    .A2(_1781_),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4364_ (.A1(_1735_),
    .A2(_1778_),
    .B(_1788_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4365_ (.I(_1364_),
    .Z(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4366_ (.I(_1777_),
    .Z(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4367_ (.I(_1780_),
    .Z(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4368_ (.A1(_1738_),
    .A2(_1791_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4369_ (.A1(_1789_),
    .A2(_1790_),
    .B(_1792_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4370_ (.A1(_1742_),
    .A2(_1791_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4371_ (.A1(_1741_),
    .A2(_1790_),
    .B(_1793_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4372_ (.A1(_1745_),
    .A2(_1791_),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4373_ (.A1(_1744_),
    .A2(_1790_),
    .B(_1794_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4374_ (.A1(_1748_),
    .A2(_1791_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4375_ (.A1(_1747_),
    .A2(_1790_),
    .B(_1795_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4376_ (.I(_1777_),
    .Z(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4377_ (.I(_1780_),
    .Z(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4378_ (.A1(_1752_),
    .A2(_1797_),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4379_ (.A1(_1750_),
    .A2(_1796_),
    .B(_1798_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4380_ (.A1(_1756_),
    .A2(_1797_),
    .ZN(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4381_ (.A1(_1755_),
    .A2(_1796_),
    .B(_1799_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4382_ (.I(net19),
    .Z(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4383_ (.A1(_1800_),
    .A2(_1797_),
    .ZN(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4384_ (.A1(_1758_),
    .A2(_1796_),
    .B(_1801_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4385_ (.I(_1378_),
    .Z(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4386_ (.A1(_1760_),
    .A2(_1797_),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4387_ (.A1(_1802_),
    .A2(_1796_),
    .B(_1803_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4388_ (.I(_1777_),
    .Z(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4389_ (.I(_1780_),
    .Z(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4390_ (.A1(_1764_),
    .A2(_1805_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4391_ (.A1(_1762_),
    .A2(_1804_),
    .B(_1806_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4392_ (.A1(_1768_),
    .A2(_1805_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4393_ (.A1(_1767_),
    .A2(_1804_),
    .B(_1807_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4394_ (.A1(_1771_),
    .A2(_1805_),
    .ZN(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4395_ (.A1(_1770_),
    .A2(_1804_),
    .B(_1808_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4396_ (.A1(_1774_),
    .A2(_1805_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4397_ (.A1(_1773_),
    .A2(_1804_),
    .B(_1809_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4398_ (.A1(_1724_),
    .A2(_1226_),
    .ZN(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4399_ (.I(_1810_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4400_ (.I(_1811_),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4401_ (.I(_1810_),
    .Z(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4402_ (.I(_1813_),
    .Z(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4403_ (.A1(_1779_),
    .A2(_1814_),
    .ZN(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4404_ (.A1(_1723_),
    .A2(_1812_),
    .B(_1815_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4405_ (.A1(_1783_),
    .A2(_1814_),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4406_ (.A1(_1731_),
    .A2(_1812_),
    .B(_1816_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4407_ (.A1(_1785_),
    .A2(_1814_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4408_ (.A1(_1733_),
    .A2(_1812_),
    .B(_1817_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4409_ (.A1(_1787_),
    .A2(_1814_),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4410_ (.A1(_1735_),
    .A2(_1812_),
    .B(_1818_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4411_ (.I(_1811_),
    .Z(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4412_ (.I(_1813_),
    .Z(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4413_ (.A1(_1738_),
    .A2(_1820_),
    .ZN(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4414_ (.A1(_1789_),
    .A2(_1819_),
    .B(_1821_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4415_ (.A1(_1742_),
    .A2(_1820_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4416_ (.A1(_1741_),
    .A2(_1819_),
    .B(_1822_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4417_ (.A1(_1745_),
    .A2(_1820_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4418_ (.A1(_1744_),
    .A2(_1819_),
    .B(_1823_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4419_ (.A1(_1748_),
    .A2(_1820_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4420_ (.A1(_1747_),
    .A2(_1819_),
    .B(_1824_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4421_ (.I(_1811_),
    .Z(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4422_ (.I(_1813_),
    .Z(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4423_ (.A1(_1752_),
    .A2(_1826_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4424_ (.A1(_1750_),
    .A2(_1825_),
    .B(_1827_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4425_ (.A1(_1756_),
    .A2(_1826_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4426_ (.A1(_1755_),
    .A2(_1825_),
    .B(_1828_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4427_ (.A1(_1800_),
    .A2(_1826_),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4428_ (.A1(_1758_),
    .A2(_1825_),
    .B(_1829_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4429_ (.A1(_1760_),
    .A2(_1826_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4430_ (.A1(_1802_),
    .A2(_1825_),
    .B(_1830_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4431_ (.I(_1811_),
    .Z(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4432_ (.I(_1813_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4433_ (.A1(_1764_),
    .A2(_1832_),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4434_ (.A1(_1762_),
    .A2(_1831_),
    .B(_1833_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4435_ (.A1(_1768_),
    .A2(_1832_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4436_ (.A1(_1767_),
    .A2(_1831_),
    .B(_1834_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4437_ (.A1(_1771_),
    .A2(_1832_),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4438_ (.A1(_1770_),
    .A2(_1831_),
    .B(_1835_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4439_ (.A1(_1774_),
    .A2(_1832_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4440_ (.A1(_1773_),
    .A2(_1831_),
    .B(_1836_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4441_ (.A1(_0931_),
    .A2(_0966_),
    .ZN(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4442_ (.I(_1837_),
    .Z(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4443_ (.I(_1838_),
    .Z(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4444_ (.I(_1837_),
    .Z(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4445_ (.I(_1840_),
    .Z(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4446_ (.A1(_1779_),
    .A2(_1841_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4447_ (.A1(_1723_),
    .A2(_1839_),
    .B(_1842_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4448_ (.A1(_1783_),
    .A2(_1841_),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4449_ (.A1(_1731_),
    .A2(_1839_),
    .B(_1843_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4450_ (.A1(_1785_),
    .A2(_1841_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4451_ (.A1(_1733_),
    .A2(_1839_),
    .B(_1844_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4452_ (.A1(_1787_),
    .A2(_1841_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4453_ (.A1(_1735_),
    .A2(_1839_),
    .B(_1845_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4454_ (.I(_1838_),
    .Z(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4455_ (.I(_1840_),
    .Z(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4456_ (.A1(_1738_),
    .A2(_1847_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4457_ (.A1(_1789_),
    .A2(_1846_),
    .B(_1848_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4458_ (.A1(_1742_),
    .A2(_1847_),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4459_ (.A1(_1741_),
    .A2(_1846_),
    .B(_1849_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4460_ (.A1(_1745_),
    .A2(_1847_),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4461_ (.A1(_1744_),
    .A2(_1846_),
    .B(_1850_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4462_ (.A1(_1748_),
    .A2(_1847_),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4463_ (.A1(_1747_),
    .A2(_1846_),
    .B(_1851_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4464_ (.I(_1838_),
    .Z(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4465_ (.I(_1840_),
    .Z(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4466_ (.A1(_1752_),
    .A2(_1853_),
    .ZN(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4467_ (.A1(_1750_),
    .A2(_1852_),
    .B(_1854_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4468_ (.A1(_1756_),
    .A2(_1853_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4469_ (.A1(_1755_),
    .A2(_1852_),
    .B(_1855_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4470_ (.A1(_1800_),
    .A2(_1853_),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4471_ (.A1(_1758_),
    .A2(_1852_),
    .B(_1856_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4472_ (.A1(_1760_),
    .A2(_1853_),
    .ZN(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4473_ (.A1(_1802_),
    .A2(_1852_),
    .B(_1857_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4474_ (.I(_1838_),
    .Z(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4475_ (.I(_1840_),
    .Z(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4476_ (.A1(_1764_),
    .A2(_1859_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4477_ (.A1(_1762_),
    .A2(_1858_),
    .B(_1860_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4478_ (.A1(_1768_),
    .A2(_1859_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4479_ (.A1(_1767_),
    .A2(_1858_),
    .B(_1861_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4480_ (.A1(_1771_),
    .A2(_1859_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4481_ (.A1(_1770_),
    .A2(_1858_),
    .B(_1862_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4482_ (.A1(_1774_),
    .A2(_1859_),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4483_ (.A1(_1773_),
    .A2(_1858_),
    .B(_1863_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4484_ (.I(_2145_),
    .Z(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4485_ (.A1(_1724_),
    .A2(_1286_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4486_ (.I(_1865_),
    .Z(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4487_ (.I(_1866_),
    .Z(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4488_ (.I(_1865_),
    .Z(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4489_ (.I(_1868_),
    .Z(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4490_ (.A1(_1779_),
    .A2(_1869_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4491_ (.A1(_1864_),
    .A2(_1867_),
    .B(_1870_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4492_ (.I(_2171_),
    .Z(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4493_ (.A1(_1783_),
    .A2(_1869_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4494_ (.A1(_1871_),
    .A2(_1867_),
    .B(_1872_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4495_ (.I(_2189_),
    .Z(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4496_ (.A1(_1785_),
    .A2(_1869_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4497_ (.A1(_1873_),
    .A2(_1867_),
    .B(_1874_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4498_ (.I(_2211_),
    .Z(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4499_ (.A1(_1787_),
    .A2(_1869_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4500_ (.A1(_1875_),
    .A2(_1867_),
    .B(_1876_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4501_ (.I(_1866_),
    .Z(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4502_ (.I(net28),
    .Z(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4503_ (.I(_1868_),
    .Z(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4504_ (.A1(_1878_),
    .A2(_1879_),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4505_ (.A1(_1789_),
    .A2(_1877_),
    .B(_1880_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4506_ (.I(_2256_),
    .Z(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4507_ (.I(net29),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4508_ (.A1(_1882_),
    .A2(_1879_),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4509_ (.A1(_1881_),
    .A2(_1877_),
    .B(_1883_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4510_ (.I(_2277_),
    .Z(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4511_ (.I(net30),
    .Z(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4512_ (.A1(_1885_),
    .A2(_1879_),
    .ZN(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4513_ (.A1(_1884_),
    .A2(_1877_),
    .B(_1886_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4514_ (.I(_2297_),
    .Z(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4515_ (.I(net31),
    .Z(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4516_ (.A1(_1888_),
    .A2(_1879_),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4517_ (.A1(_1887_),
    .A2(_1877_),
    .B(_1889_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4518_ (.I(_2321_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4519_ (.I(_1866_),
    .Z(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4520_ (.I(net32),
    .Z(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4521_ (.I(_1868_),
    .Z(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4522_ (.A1(_1892_),
    .A2(_1893_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4523_ (.A1(_1890_),
    .A2(_1891_),
    .B(_1894_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4524_ (.I(_2335_),
    .Z(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4525_ (.I(net33),
    .Z(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4526_ (.A1(_1896_),
    .A2(_1893_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4527_ (.A1(_1895_),
    .A2(_1891_),
    .B(_1897_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4528_ (.I(_2354_),
    .Z(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4529_ (.A1(_1800_),
    .A2(_1893_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4530_ (.A1(_1898_),
    .A2(_1891_),
    .B(_1899_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4531_ (.I(net20),
    .Z(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4532_ (.A1(_1900_),
    .A2(_1893_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4533_ (.A1(_1802_),
    .A2(_1891_),
    .B(_1901_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4534_ (.I(_0571_),
    .Z(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4535_ (.I(_1866_),
    .Z(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4536_ (.I(net21),
    .Z(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4537_ (.I(_1868_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4538_ (.A1(_1904_),
    .A2(_1905_),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4539_ (.A1(_1902_),
    .A2(_1903_),
    .B(_1906_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4540_ (.I(_0591_),
    .Z(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4541_ (.I(net22),
    .Z(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4542_ (.A1(_1908_),
    .A2(_1905_),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4543_ (.A1(_1907_),
    .A2(_1903_),
    .B(_1909_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4544_ (.I(_0603_),
    .Z(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4545_ (.I(net23),
    .Z(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4546_ (.A1(_1911_),
    .A2(_1905_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4547_ (.A1(_1910_),
    .A2(_1903_),
    .B(_1912_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4548_ (.I(_0614_),
    .Z(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4549_ (.I(net24),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4550_ (.A1(_1914_),
    .A2(_1905_),
    .ZN(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4551_ (.A1(_1913_),
    .A2(_1903_),
    .B(_1915_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4552_ (.A1(_1724_),
    .A2(_1033_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4553_ (.I(_1916_),
    .Z(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4554_ (.I(_1917_),
    .Z(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4555_ (.I(net18),
    .Z(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4556_ (.I(_1916_),
    .Z(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4557_ (.I(_1920_),
    .Z(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4558_ (.A1(_1919_),
    .A2(_1921_),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4559_ (.A1(_1864_),
    .A2(_1918_),
    .B(_1922_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4560_ (.I(net25),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4561_ (.A1(_1923_),
    .A2(_1921_),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4562_ (.A1(_1871_),
    .A2(_1918_),
    .B(_1924_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4563_ (.I(net26),
    .Z(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4564_ (.A1(_1925_),
    .A2(_1921_),
    .ZN(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4565_ (.A1(_1873_),
    .A2(_1918_),
    .B(_1926_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4566_ (.I(net27),
    .Z(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4567_ (.A1(_1927_),
    .A2(_1921_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4568_ (.A1(_1875_),
    .A2(_1918_),
    .B(_1928_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4569_ (.I(_2232_),
    .Z(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4570_ (.I(_1917_),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4571_ (.I(_1920_),
    .Z(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4572_ (.A1(_1878_),
    .A2(_1931_),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4573_ (.A1(_1929_),
    .A2(_1930_),
    .B(_1932_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4574_ (.A1(_1882_),
    .A2(_1931_),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4575_ (.A1(_1881_),
    .A2(_1930_),
    .B(_1933_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4576_ (.A1(_1885_),
    .A2(_1931_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4577_ (.A1(_1884_),
    .A2(_1930_),
    .B(_1934_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4578_ (.A1(_1888_),
    .A2(_1931_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4579_ (.A1(_1887_),
    .A2(_1930_),
    .B(_1935_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4580_ (.I(_1917_),
    .Z(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4581_ (.I(_1920_),
    .Z(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4582_ (.A1(_1892_),
    .A2(_1937_),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4583_ (.A1(_1890_),
    .A2(_1936_),
    .B(_1938_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4584_ (.A1(_1896_),
    .A2(_1937_),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4585_ (.A1(_1895_),
    .A2(_1936_),
    .B(_1939_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4586_ (.I(net19),
    .Z(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4587_ (.A1(_1940_),
    .A2(_1937_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4588_ (.A1(_1898_),
    .A2(_1936_),
    .B(_1941_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4589_ (.I(_2370_),
    .Z(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4590_ (.A1(_1900_),
    .A2(_1937_),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4591_ (.A1(_1942_),
    .A2(_1936_),
    .B(_1943_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4592_ (.I(_1917_),
    .Z(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4593_ (.I(_1920_),
    .Z(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4594_ (.A1(_1904_),
    .A2(_1945_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4595_ (.A1(_1902_),
    .A2(_1944_),
    .B(_1946_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4596_ (.A1(_1908_),
    .A2(_1945_),
    .ZN(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4597_ (.A1(_1907_),
    .A2(_1944_),
    .B(_1947_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4598_ (.A1(_1911_),
    .A2(_1945_),
    .ZN(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4599_ (.A1(_1910_),
    .A2(_1944_),
    .B(_1948_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4600_ (.A1(_1914_),
    .A2(_1945_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4601_ (.A1(_1913_),
    .A2(_1944_),
    .B(_1949_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4602_ (.A1(_0966_),
    .A2(_1068_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4603_ (.I(_1950_),
    .Z(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4604_ (.I(_1951_),
    .Z(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4605_ (.I(_1950_),
    .Z(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4606_ (.I(_1953_),
    .Z(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4607_ (.A1(_1919_),
    .A2(_1954_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4608_ (.A1(_1864_),
    .A2(_1952_),
    .B(_1955_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4609_ (.A1(_1923_),
    .A2(_1954_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4610_ (.A1(_1871_),
    .A2(_1952_),
    .B(_1956_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4611_ (.A1(_1925_),
    .A2(_1954_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4612_ (.A1(_1873_),
    .A2(_1952_),
    .B(_1957_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4613_ (.A1(_1927_),
    .A2(_1954_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4614_ (.A1(_1875_),
    .A2(_1952_),
    .B(_1958_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4615_ (.I(_1951_),
    .Z(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4616_ (.I(_1953_),
    .Z(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4617_ (.A1(_1878_),
    .A2(_1960_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4618_ (.A1(_1929_),
    .A2(_1959_),
    .B(_1961_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4619_ (.A1(_1882_),
    .A2(_1960_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4620_ (.A1(_1881_),
    .A2(_1959_),
    .B(_1962_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4621_ (.A1(_1885_),
    .A2(_1960_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4622_ (.A1(_1884_),
    .A2(_1959_),
    .B(_1963_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4623_ (.A1(_1888_),
    .A2(_1960_),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4624_ (.A1(_1887_),
    .A2(_1959_),
    .B(_1964_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4625_ (.I(_1951_),
    .Z(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4626_ (.I(_1953_),
    .Z(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4627_ (.A1(_1892_),
    .A2(_1966_),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4628_ (.A1(_1890_),
    .A2(_1965_),
    .B(_1967_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4629_ (.A1(_1896_),
    .A2(_1966_),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4630_ (.A1(_1895_),
    .A2(_1965_),
    .B(_1968_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4631_ (.A1(_1940_),
    .A2(_1966_),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4632_ (.A1(_1898_),
    .A2(_1965_),
    .B(_1969_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4633_ (.A1(_1900_),
    .A2(_1966_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4634_ (.A1(_1942_),
    .A2(_1965_),
    .B(_1970_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4635_ (.I(_1951_),
    .Z(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4636_ (.I(_1953_),
    .Z(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4637_ (.A1(_1904_),
    .A2(_1972_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4638_ (.A1(_1902_),
    .A2(_1971_),
    .B(_1973_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4639_ (.A1(_1908_),
    .A2(_1972_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4640_ (.A1(_1907_),
    .A2(_1971_),
    .B(_1974_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4641_ (.A1(_1911_),
    .A2(_1972_),
    .ZN(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4642_ (.A1(_1910_),
    .A2(_1971_),
    .B(_1975_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4643_ (.A1(_1914_),
    .A2(_1972_),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4644_ (.A1(_1913_),
    .A2(_1971_),
    .B(_1976_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4645_ (.A1(_0933_),
    .A2(_1226_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4646_ (.I(_1977_),
    .Z(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4647_ (.I(_1978_),
    .Z(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4648_ (.I(_1977_),
    .Z(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4649_ (.I(_1980_),
    .Z(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4650_ (.A1(_1919_),
    .A2(_1981_),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4651_ (.A1(_1864_),
    .A2(_1979_),
    .B(_1982_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4652_ (.A1(_1923_),
    .A2(_1981_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4653_ (.A1(_1871_),
    .A2(_1979_),
    .B(_1983_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4654_ (.A1(_1925_),
    .A2(_1981_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4655_ (.A1(_1873_),
    .A2(_1979_),
    .B(_1984_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4656_ (.A1(_1927_),
    .A2(_1981_),
    .ZN(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4657_ (.A1(_1875_),
    .A2(_1979_),
    .B(_1985_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4658_ (.I(_1978_),
    .Z(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4659_ (.I(_1980_),
    .Z(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4660_ (.A1(_1878_),
    .A2(_1987_),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4661_ (.A1(_1929_),
    .A2(_1986_),
    .B(_1988_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4662_ (.A1(_1882_),
    .A2(_1987_),
    .ZN(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4663_ (.A1(_1881_),
    .A2(_1986_),
    .B(_1989_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4664_ (.A1(_1885_),
    .A2(_1987_),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4665_ (.A1(_1884_),
    .A2(_1986_),
    .B(_1990_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4666_ (.A1(_1888_),
    .A2(_1987_),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4667_ (.A1(_1887_),
    .A2(_1986_),
    .B(_1991_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4668_ (.I(_1978_),
    .Z(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4669_ (.I(_1980_),
    .Z(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4670_ (.A1(_1892_),
    .A2(_1993_),
    .ZN(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4671_ (.A1(_1890_),
    .A2(_1992_),
    .B(_1994_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4672_ (.A1(_1896_),
    .A2(_1993_),
    .ZN(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4673_ (.A1(_1895_),
    .A2(_1992_),
    .B(_1995_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4674_ (.A1(_1940_),
    .A2(_1993_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4675_ (.A1(_1898_),
    .A2(_1992_),
    .B(_1996_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4676_ (.A1(_1900_),
    .A2(_1993_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4677_ (.A1(_1942_),
    .A2(_1992_),
    .B(_1997_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4678_ (.I(_1978_),
    .Z(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4679_ (.I(_1980_),
    .Z(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4680_ (.A1(_1904_),
    .A2(_1999_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4681_ (.A1(_1902_),
    .A2(_1998_),
    .B(_2000_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4682_ (.A1(_1908_),
    .A2(_1999_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4683_ (.A1(_1907_),
    .A2(_1998_),
    .B(_2001_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4684_ (.A1(_1911_),
    .A2(_1999_),
    .ZN(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4685_ (.A1(_1910_),
    .A2(_1998_),
    .B(_2002_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4686_ (.A1(_1914_),
    .A2(_1999_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4687_ (.A1(_1913_),
    .A2(_1998_),
    .B(_2003_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4688_ (.A1(_0933_),
    .A2(_1286_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4689_ (.I(_2004_),
    .Z(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4690_ (.I(_2005_),
    .Z(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4691_ (.I(_2004_),
    .Z(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4692_ (.I(_2007_),
    .Z(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4693_ (.A1(_1919_),
    .A2(_2008_),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4694_ (.A1(_0961_),
    .A2(_2006_),
    .B(_2009_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4695_ (.A1(_1923_),
    .A2(_2008_),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4696_ (.A1(_0973_),
    .A2(_2006_),
    .B(_2010_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4697_ (.A1(_1925_),
    .A2(_2008_),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4698_ (.A1(_0976_),
    .A2(_2006_),
    .B(_2011_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4699_ (.A1(_1927_),
    .A2(_2008_),
    .ZN(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4700_ (.A1(_0979_),
    .A2(_2006_),
    .B(_2012_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4701_ (.I(_2005_),
    .Z(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4702_ (.I(_2007_),
    .Z(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4703_ (.A1(_0797_),
    .A2(_2014_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4704_ (.A1(_1929_),
    .A2(_2013_),
    .B(_2015_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4705_ (.A1(_0801_),
    .A2(_2014_),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4706_ (.A1(_0986_),
    .A2(_2013_),
    .B(_2016_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4707_ (.A1(_0804_),
    .A2(_2014_),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4708_ (.A1(_0990_),
    .A2(_2013_),
    .B(_2017_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4709_ (.A1(_0807_),
    .A2(_2014_),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4710_ (.A1(_0994_),
    .A2(_2013_),
    .B(_2018_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4711_ (.I(_2005_),
    .Z(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4712_ (.I(_2007_),
    .Z(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4713_ (.A1(_0811_),
    .A2(_2020_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4714_ (.A1(_0998_),
    .A2(_2019_),
    .B(_2021_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4715_ (.A1(_0815_),
    .A2(_2020_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4716_ (.A1(_1004_),
    .A2(_2019_),
    .B(_2022_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4717_ (.A1(_1940_),
    .A2(_2020_),
    .ZN(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4718_ (.A1(_1008_),
    .A2(_2019_),
    .B(_2023_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4719_ (.A1(_0823_),
    .A2(_2020_),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4720_ (.A1(_1942_),
    .A2(_2019_),
    .B(_2024_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4721_ (.I(_2005_),
    .Z(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4722_ (.I(_2007_),
    .Z(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4723_ (.A1(_0827_),
    .A2(_2026_),
    .ZN(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4724_ (.A1(_1013_),
    .A2(_2025_),
    .B(_2027_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4725_ (.A1(_0831_),
    .A2(_2026_),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4726_ (.A1(_1019_),
    .A2(_2025_),
    .B(_2028_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4727_ (.A1(_0834_),
    .A2(_2026_),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4728_ (.A1(_1023_),
    .A2(_2025_),
    .B(_2029_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4729_ (.A1(_0837_),
    .A2(_2026_),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4730_ (.A1(_1027_),
    .A2(_2025_),
    .B(_2030_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4731_ (.A1(_1068_),
    .A2(_1414_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4732_ (.I(_2031_),
    .Z(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4733_ (.I(_2032_),
    .Z(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4734_ (.I(_2031_),
    .Z(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4735_ (.I(_2034_),
    .Z(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4736_ (.A1(_0780_),
    .A2(_2035_),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4737_ (.A1(_0961_),
    .A2(_2033_),
    .B(_2036_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4738_ (.A1(_0785_),
    .A2(_2035_),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4739_ (.A1(_0973_),
    .A2(_2033_),
    .B(_2037_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4740_ (.A1(_0788_),
    .A2(_2035_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4741_ (.A1(_0976_),
    .A2(_2033_),
    .B(_2038_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4742_ (.A1(_0791_),
    .A2(_2035_),
    .ZN(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4743_ (.A1(_0979_),
    .A2(_2033_),
    .B(_2039_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4744_ (.I(_2032_),
    .Z(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4745_ (.I(_2034_),
    .Z(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4746_ (.A1(_0797_),
    .A2(_2041_),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4747_ (.A1(_0794_),
    .A2(_2040_),
    .B(_2042_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4748_ (.A1(_0801_),
    .A2(_2041_),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4749_ (.A1(_0986_),
    .A2(_2040_),
    .B(_2043_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4750_ (.A1(_0804_),
    .A2(_2041_),
    .ZN(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4751_ (.A1(_0990_),
    .A2(_2040_),
    .B(_2044_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4752_ (.A1(_0807_),
    .A2(_2041_),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4753_ (.A1(_0994_),
    .A2(_2040_),
    .B(_2045_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4754_ (.I(_2032_),
    .Z(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4755_ (.I(_2034_),
    .Z(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4756_ (.A1(_0811_),
    .A2(_2047_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4757_ (.A1(_0998_),
    .A2(_2046_),
    .B(_2048_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4758_ (.A1(_0815_),
    .A2(_2047_),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4759_ (.A1(_1004_),
    .A2(_2046_),
    .B(_2049_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4760_ (.A1(_0818_),
    .A2(_2047_),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4761_ (.A1(_1008_),
    .A2(_2046_),
    .B(_2050_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4762_ (.A1(_0823_),
    .A2(_2047_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4763_ (.A1(_0821_),
    .A2(_2046_),
    .B(_2051_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4764_ (.I(_2032_),
    .Z(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4765_ (.I(_2034_),
    .Z(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4766_ (.A1(_0827_),
    .A2(_2053_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4767_ (.A1(_1013_),
    .A2(_2052_),
    .B(_2054_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4768_ (.A1(_0831_),
    .A2(_2053_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4769_ (.A1(_1019_),
    .A2(_2052_),
    .B(_2055_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4770_ (.A1(_0834_),
    .A2(_2053_),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4771_ (.A1(_1023_),
    .A2(_2052_),
    .B(_2056_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4772_ (.A1(_0837_),
    .A2(_2053_),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4773_ (.A1(_1027_),
    .A2(_2052_),
    .B(_2057_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4774_ (.I(net47),
    .Z(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4775_ (.A1(_2058_),
    .A2(_0731_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4776_ (.A1(_2145_),
    .A2(_0752_),
    .B1(_0713_),
    .B2(_2119_),
    .ZN(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4777_ (.A1(net35),
    .A2(_2059_),
    .A3(_2060_),
    .ZN(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4778_ (.A1(_0718_),
    .A2(_2061_),
    .Z(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4779_ (.I(_2062_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4780_ (.I(net51),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4781_ (.A1(_2058_),
    .A2(_2063_),
    .Z(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4782_ (.A1(_2171_),
    .A2(_0753_),
    .B1(_0732_),
    .B2(_2064_),
    .C(_0708_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4783_ (.A1(_2084_),
    .A2(_0667_),
    .B(_2065_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4784_ (.A1(_2063_),
    .A2(_0730_),
    .B(_2066_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4785_ (.I(net52),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4786_ (.A1(_2058_),
    .A2(net51),
    .A3(net52),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4787_ (.A1(_2058_),
    .A2(net51),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4788_ (.A1(_2067_),
    .A2(_2069_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4789_ (.A1(_2068_),
    .A2(_2070_),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4790_ (.A1(_2189_),
    .A2(_0753_),
    .B1(_0732_),
    .B2(_2071_),
    .C(_0708_),
    .ZN(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4791_ (.A1(_0688_),
    .A2(_0667_),
    .B(_2072_),
    .ZN(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4792_ (.A1(_2067_),
    .A2(_0730_),
    .B(_2073_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4793_ (.A1(_2211_),
    .A2(_0753_),
    .Z(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4794_ (.I(net53),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4795_ (.A1(_2075_),
    .A2(_2068_),
    .Z(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4796_ (.A1(\Control_unit2.instr_stage2[3] ),
    .A2(_0747_),
    .B1(_0713_),
    .B2(_2076_),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4797_ (.A1(_0709_),
    .A2(_2074_),
    .A3(_2077_),
    .B1(_0749_),
    .B2(_2075_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4798_ (.D(_0000_),
    .RN(net34),
    .CLK(clknet_leaf_7_clk),
    .Q(net54));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4799_ (.D(_0001_),
    .RN(net34),
    .CLK(clknet_leaf_6_clk),
    .Q(net55));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4800_ (.D(_0002_),
    .RN(net34),
    .CLK(clknet_leaf_14_clk),
    .Q(net56));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4801_ (.D(_0003_),
    .RN(net34),
    .CLK(clknet_leaf_6_clk),
    .Q(net57));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4802_ (.D(_0004_),
    .RN(net34),
    .CLK(clknet_leaf_6_clk),
    .Q(net58));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4803_ (.D(_0005_),
    .RN(net34),
    .CLK(clknet_leaf_11_clk),
    .Q(net59));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4804_ (.D(_0006_),
    .RN(net34),
    .CLK(clknet_leaf_6_clk),
    .Q(net48));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4805_ (.D(_0007_),
    .RN(net34),
    .CLK(clknet_leaf_15_clk),
    .Q(net49));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4806_ (.D(_0008_),
    .RN(net34),
    .CLK(clknet_leaf_15_clk),
    .Q(net50));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4807_ (.D(_0009_),
    .RN(net34),
    .CLK(clknet_leaf_34_clk),
    .Q(net60));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4808_ (.D(_0010_),
    .RN(net34),
    .CLK(clknet_leaf_33_clk),
    .Q(net67));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4809_ (.D(_0011_),
    .RN(net34),
    .CLK(clknet_leaf_34_clk),
    .Q(net68));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4810_ (.D(_0012_),
    .RN(net34),
    .CLK(clknet_leaf_34_clk),
    .Q(net69));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4811_ (.D(_0013_),
    .RN(net34),
    .CLK(clknet_leaf_37_clk),
    .Q(net70));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4812_ (.D(_0014_),
    .RN(net34),
    .CLK(clknet_leaf_36_clk),
    .Q(net71));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4813_ (.D(_0015_),
    .RN(net34),
    .CLK(clknet_leaf_36_clk),
    .Q(net72));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4814_ (.D(_0016_),
    .RN(net34),
    .CLK(clknet_leaf_36_clk),
    .Q(net73));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4815_ (.D(_0017_),
    .RN(net34),
    .CLK(clknet_leaf_42_clk),
    .Q(net74));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4816_ (.D(_0018_),
    .RN(net34),
    .CLK(clknet_leaf_42_clk),
    .Q(net75));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4817_ (.D(_0019_),
    .RN(net34),
    .CLK(clknet_leaf_42_clk),
    .Q(net61));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4818_ (.D(_0020_),
    .RN(net34),
    .CLK(clknet_leaf_42_clk),
    .Q(net62));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4819_ (.D(_0021_),
    .RN(net34),
    .CLK(clknet_leaf_42_clk),
    .Q(net63));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4820_ (.D(_0022_),
    .RN(net34),
    .CLK(clknet_leaf_44_clk),
    .Q(net64));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4821_ (.D(_0023_),
    .RN(net34),
    .CLK(clknet_leaf_44_clk),
    .Q(net65));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4822_ (.D(_0024_),
    .RN(net34),
    .CLK(clknet_leaf_44_clk),
    .Q(net66));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4823_ (.D(_0025_),
    .RN(net34),
    .CLK(clknet_leaf_4_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[0].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4824_ (.D(_0026_),
    .RN(net34),
    .CLK(clknet_leaf_21_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[1].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4825_ (.D(_0027_),
    .RN(net34),
    .CLK(clknet_leaf_21_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[2].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4826_ (.D(_0028_),
    .RN(net34),
    .CLK(clknet_leaf_15_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[3].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4827_ (.D(_0029_),
    .RN(net34),
    .CLK(clknet_leaf_15_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[4].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4828_ (.D(_0030_),
    .RN(net34),
    .CLK(clknet_leaf_15_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4829_ (.D(_0031_),
    .RN(net34),
    .CLK(clknet_leaf_19_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[6].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4830_ (.D(_0032_),
    .RN(net34),
    .CLK(clknet_leaf_19_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[7].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4831_ (.D(_0033_),
    .RN(net34),
    .CLK(clknet_leaf_19_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4832_ (.D(_0034_),
    .RN(net34),
    .CLK(clknet_leaf_19_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i0 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4833_ (.D(_0035_),
    .RN(net34),
    .CLK(clknet_4_6_0_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4834_ (.D(_0036_),
    .RN(net34),
    .CLK(clknet_leaf_31_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[11].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4835_ (.D(_0037_),
    .RN(net34),
    .CLK(clknet_leaf_32_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[12].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4836_ (.D(_0038_),
    .RN(net34),
    .CLK(clknet_leaf_33_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[13].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4837_ (.D(_0039_),
    .RN(net34),
    .CLK(clknet_leaf_33_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[14].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4838_ (.D(_0040_),
    .RN(net34),
    .CLK(clknet_4_7_0_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.Y_CY[0].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4839_ (.D(_0041_),
    .RN(net34),
    .CLK(clknet_leaf_19_clk),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4840_ (.D(_0042_),
    .RN(net34),
    .CLK(clknet_4_7_0_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4841_ (.D(_0043_),
    .RN(net34),
    .CLK(clknet_leaf_33_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4842_ (.D(_0044_),
    .RN(net34),
    .CLK(clknet_leaf_33_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4843_ (.D(_0045_),
    .RN(net34),
    .CLK(clknet_leaf_34_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4844_ (.D(_0046_),
    .RN(net34),
    .CLK(clknet_leaf_37_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4845_ (.D(_0047_),
    .RN(net34),
    .CLK(clknet_leaf_36_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4846_ (.D(_0048_),
    .RN(net34),
    .CLK(clknet_leaf_36_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4847_ (.D(_0049_),
    .RN(net34),
    .CLK(clknet_leaf_37_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4848_ (.D(_0050_),
    .RN(net34),
    .CLK(clknet_leaf_42_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4849_ (.D(_0051_),
    .RN(net34),
    .CLK(clknet_leaf_42_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4850_ (.D(_0052_),
    .RN(net34),
    .CLK(clknet_leaf_41_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4851_ (.D(_0053_),
    .RN(net34),
    .CLK(clknet_leaf_41_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4852_ (.D(_0054_),
    .RN(net34),
    .CLK(clknet_leaf_43_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4853_ (.D(_0055_),
    .RN(net34),
    .CLK(clknet_leaf_44_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4854_ (.D(_0056_),
    .RN(net34),
    .CLK(clknet_leaf_45_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4855_ (.D(_0057_),
    .RN(net34),
    .CLK(clknet_leaf_45_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4856_ (.D(\Stack_pointer.SP_next[0] ),
    .RN(net34),
    .CLK(clknet_4_5_0_clk),
    .Q(\Stack_pointer.SP[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4857_ (.D(\Stack_pointer.SP_next[1] ),
    .RN(net34),
    .CLK(clknet_leaf_10_clk),
    .Q(\Stack_pointer.SP[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4858_ (.D(\Stack_pointer.SP_next[2] ),
    .RN(net34),
    .CLK(clknet_leaf_8_clk),
    .Q(\Stack_pointer.SP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4859_ (.D(\Stack_pointer.SP_next[3] ),
    .RN(net34),
    .CLK(clknet_leaf_8_clk),
    .Q(\Stack_pointer.SP[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _4860_ (.D(\Stack_pointer.SP_next[4] ),
    .SETN(net34),
    .CLK(clknet_leaf_10_clk),
    .Q(\Stack_pointer.SP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _4861_ (.D(\Stack_pointer.SP_next[5] ),
    .SETN(net34),
    .CLK(clknet_leaf_11_clk),
    .Q(\Stack_pointer.SP[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _4862_ (.D(\Stack_pointer.SP_next[6] ),
    .SETN(net34),
    .CLK(clknet_leaf_11_clk),
    .Q(\Stack_pointer.SP[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffsnq_1 _4863_ (.D(\Stack_pointer.SP_next[7] ),
    .SETN(net34),
    .CLK(clknet_leaf_11_clk),
    .Q(\Stack_pointer.SP[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4864_ (.D(_0058_),
    .RN(net34),
    .CLK(clknet_leaf_19_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_001.p_Z ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4865_ (.D(\Control_unit1.instr_stage1[0] ),
    .RN(net34),
    .CLK(clknet_leaf_17_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_000.ALU_func[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4866_ (.D(\Control_unit1.instr_stage1[1] ),
    .RN(net34),
    .CLK(clknet_leaf_17_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_000.ALU_func[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4867_ (.D(\Control_unit1.instr_stage1[2] ),
    .RN(net34),
    .CLK(clknet_leaf_17_clk),
    .Q(\Arithmetic_Logic_Unit.ALU_000.ALU_func[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4868_ (.D(\Control_unit1.instr_stage1[3] ),
    .RN(net34),
    .CLK(clknet_leaf_12_clk),
    .Q(\Control_unit2.instr_stage2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4869_ (.D(\Control_unit1.instr_stage1[4] ),
    .RN(net34),
    .CLK(clknet_leaf_13_clk),
    .Q(\Control_unit2.instr_stage2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4870_ (.D(\Control_unit1.instr_stage1[5] ),
    .RN(net34),
    .CLK(clknet_leaf_12_clk),
    .Q(\Control_unit2.instr_stage2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4871_ (.D(\Control_unit1.instr_stage1[6] ),
    .RN(net34),
    .CLK(clknet_leaf_13_clk),
    .Q(\Control_unit2.instr_stage2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4872_ (.D(\Control_unit1.instr_stage1[7] ),
    .RN(net34),
    .CLK(clknet_leaf_13_clk),
    .Q(\Control_unit2.instr_stage2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4873_ (.D(\Control_unit1.instr_stage1[8] ),
    .RN(net34),
    .CLK(clknet_leaf_5_clk),
    .Q(\Control_unit2.instr_stage2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4874_ (.D(\Control_unit1.instr_stage1[9] ),
    .RN(net34),
    .CLK(clknet_leaf_5_clk),
    .Q(\Control_unit2.instr_stage2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4875_ (.D(\Control_unit1.instr_stage1[10] ),
    .RN(net34),
    .CLK(clknet_leaf_4_clk),
    .Q(\Control_unit2.instr_stage2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4876_ (.D(\Control_unit1.instr_stage1[11] ),
    .RN(net34),
    .CLK(clknet_leaf_17_clk),
    .Q(\Control_unit2.instr_stage2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4877_ (.D(\Control_unit1.instr_stage1[12] ),
    .RN(net34),
    .CLK(clknet_leaf_4_clk),
    .Q(\Control_unit2.instr_stage2[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4878_ (.D(\Control_unit1.instr_decoder1.A[0] ),
    .RN(net34),
    .CLK(clknet_leaf_18_clk),
    .Q(\Arithmetic_Logic_Unit.op ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_2 _4879_ (.D(\Control_unit1.instr_decoder1.A[1] ),
    .RN(net34),
    .CLK(clknet_leaf_18_clk),
    .Q(\Control_unit2.instr_decoder2.A[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4880_ (.D(\Control_unit1.instr_decoder1.A[2] ),
    .RN(net34),
    .CLK(clknet_leaf_18_clk),
    .Q(\Control_unit2.instr_decoder2.A[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4881_ (.D(net2),
    .RN(net34),
    .CLK(clknet_leaf_8_clk),
    .Q(\Control_unit1.instr_stage1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4882_ (.D(net9),
    .RN(net34),
    .CLK(clknet_leaf_8_clk),
    .Q(\Control_unit1.instr_stage1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4883_ (.D(net10),
    .RN(net34),
    .CLK(clknet_leaf_8_clk),
    .Q(\Control_unit1.instr_stage1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4884_ (.D(net11),
    .RN(net34),
    .CLK(clknet_leaf_8_clk),
    .Q(\Control_unit1.instr_stage1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4885_ (.D(net12),
    .RN(net34),
    .CLK(clknet_leaf_8_clk),
    .Q(\Control_unit1.instr_stage1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4886_ (.D(net13),
    .RN(net34),
    .CLK(clknet_leaf_8_clk),
    .Q(\Control_unit1.instr_stage1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4887_ (.D(net14),
    .RN(net34),
    .CLK(clknet_leaf_8_clk),
    .Q(\Control_unit1.instr_stage1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4888_ (.D(net15),
    .RN(net34),
    .CLK(clknet_leaf_8_clk),
    .Q(\Control_unit1.instr_stage1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4889_ (.D(net16),
    .RN(net34),
    .CLK(clknet_leaf_7_clk),
    .Q(\Control_unit1.instr_stage1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4890_ (.D(net17),
    .RN(net34),
    .CLK(clknet_leaf_11_clk),
    .Q(\Control_unit1.instr_stage1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4891_ (.D(net3),
    .RN(net34),
    .CLK(clknet_leaf_12_clk),
    .Q(\Control_unit1.instr_stage1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4892_ (.D(net4),
    .RN(net34),
    .CLK(clknet_leaf_12_clk),
    .Q(\Control_unit1.instr_stage1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4893_ (.D(net5),
    .RN(net34),
    .CLK(clknet_leaf_12_clk),
    .Q(\Control_unit1.instr_stage1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4894_ (.D(net6),
    .RN(net34),
    .CLK(clknet_leaf_18_clk),
    .Q(\Control_unit1.instr_decoder1.A[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4895_ (.D(net7),
    .RN(net34),
    .CLK(clknet_leaf_18_clk),
    .Q(\Control_unit1.instr_decoder1.A[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4896_ (.D(net8),
    .RN(net34),
    .CLK(clknet_leaf_18_clk),
    .Q(\Control_unit1.instr_decoder1.A[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4897_ (.D(_0059_),
    .RN(net34),
    .CLK(clknet_leaf_32_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4898_ (.D(_0060_),
    .RN(net34),
    .CLK(clknet_leaf_33_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4899_ (.D(_0061_),
    .RN(net34),
    .CLK(clknet_leaf_33_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4900_ (.D(_0062_),
    .RN(net34),
    .CLK(clknet_leaf_32_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4901_ (.D(_0063_),
    .RN(net34),
    .CLK(clknet_leaf_37_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4902_ (.D(_0064_),
    .RN(net34),
    .CLK(clknet_leaf_36_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4903_ (.D(_0065_),
    .RN(net34),
    .CLK(clknet_leaf_36_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4904_ (.D(_0066_),
    .RN(net34),
    .CLK(clknet_leaf_37_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4905_ (.D(_0067_),
    .RN(net34),
    .CLK(clknet_leaf_42_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4906_ (.D(_0068_),
    .RN(net34),
    .CLK(clknet_leaf_36_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4907_ (.D(_0069_),
    .RN(net34),
    .CLK(clknet_leaf_41_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4908_ (.D(_0070_),
    .RN(net34),
    .CLK(clknet_leaf_37_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4909_ (.D(_0071_),
    .RN(net34),
    .CLK(clknet_leaf_43_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4910_ (.D(_0072_),
    .RN(net34),
    .CLK(clknet_leaf_44_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4911_ (.D(_0073_),
    .RN(net34),
    .CLK(clknet_leaf_45_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4912_ (.D(_0074_),
    .RN(net34),
    .CLK(clknet_leaf_45_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4913_ (.D(_0075_),
    .RN(net34),
    .CLK(clknet_leaf_32_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4914_ (.D(_0076_),
    .RN(net34),
    .CLK(clknet_leaf_31_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4915_ (.D(_0077_),
    .RN(net34),
    .CLK(clknet_leaf_31_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4916_ (.D(_0078_),
    .RN(net34),
    .CLK(clknet_leaf_30_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4917_ (.D(_0079_),
    .RN(net34),
    .CLK(clknet_leaf_38_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4918_ (.D(_0080_),
    .RN(net34),
    .CLK(clknet_leaf_38_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4919_ (.D(_0081_),
    .RN(net34),
    .CLK(clknet_leaf_38_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4920_ (.D(_0082_),
    .RN(net34),
    .CLK(clknet_leaf_38_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4921_ (.D(_0083_),
    .RN(net34),
    .CLK(clknet_leaf_40_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4922_ (.D(_0084_),
    .RN(net34),
    .CLK(clknet_leaf_41_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4923_ (.D(_0085_),
    .RN(net34),
    .CLK(clknet_leaf_40_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4924_ (.D(_0086_),
    .RN(net34),
    .CLK(clknet_leaf_40_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4925_ (.D(_0087_),
    .RN(net34),
    .CLK(clknet_leaf_46_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4926_ (.D(_0088_),
    .RN(net34),
    .CLK(clknet_leaf_46_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4927_ (.D(_0089_),
    .RN(net34),
    .CLK(clknet_leaf_45_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4928_ (.D(_0090_),
    .RN(net34),
    .CLK(clknet_leaf_45_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4929_ (.D(_0091_),
    .RN(net34),
    .CLK(clknet_leaf_27_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4930_ (.D(_0092_),
    .RN(net34),
    .CLK(clknet_leaf_24_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4931_ (.D(_0093_),
    .RN(net34),
    .CLK(clknet_leaf_26_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4932_ (.D(_0094_),
    .RN(net34),
    .CLK(clknet_leaf_27_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4933_ (.D(_0095_),
    .RN(net34),
    .CLK(clknet_leaf_28_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4934_ (.D(_0096_),
    .RN(net34),
    .CLK(clknet_leaf_28_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4935_ (.D(_0097_),
    .RN(net34),
    .CLK(clknet_leaf_28_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4936_ (.D(_0098_),
    .RN(net34),
    .CLK(clknet_leaf_28_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4937_ (.D(_0099_),
    .RN(net34),
    .CLK(clknet_leaf_50_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4938_ (.D(_0100_),
    .RN(net34),
    .CLK(clknet_leaf_50_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4939_ (.D(_0101_),
    .RN(net34),
    .CLK(clknet_leaf_51_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4940_ (.D(_0102_),
    .RN(net34),
    .CLK(clknet_leaf_51_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4941_ (.D(_0103_),
    .RN(net34),
    .CLK(clknet_leaf_48_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4942_ (.D(_0104_),
    .RN(net34),
    .CLK(clknet_leaf_47_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4943_ (.D(_0105_),
    .RN(net34),
    .CLK(clknet_leaf_47_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4944_ (.D(_0106_),
    .RN(net34),
    .CLK(clknet_leaf_47_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4945_ (.D(_0107_),
    .RN(net34),
    .CLK(clknet_leaf_26_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4946_ (.D(_0108_),
    .RN(net34),
    .CLK(clknet_leaf_26_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4947_ (.D(_0109_),
    .RN(net34),
    .CLK(clknet_leaf_31_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4948_ (.D(_0110_),
    .RN(net34),
    .CLK(clknet_leaf_30_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4949_ (.D(_0111_),
    .RN(net34),
    .CLK(clknet_leaf_28_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4950_ (.D(_0112_),
    .RN(net34),
    .CLK(clknet_4_13_0_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4951_ (.D(_0113_),
    .RN(net34),
    .CLK(clknet_leaf_39_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4952_ (.D(_0114_),
    .RN(net34),
    .CLK(clknet_leaf_39_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4953_ (.D(_0115_),
    .RN(net34),
    .CLK(clknet_leaf_49_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4954_ (.D(_0116_),
    .RN(net34),
    .CLK(clknet_leaf_40_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4955_ (.D(_0117_),
    .RN(net34),
    .CLK(clknet_leaf_49_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4956_ (.D(_0118_),
    .RN(net34),
    .CLK(clknet_leaf_50_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4957_ (.D(_0119_),
    .RN(net34),
    .CLK(clknet_leaf_49_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4958_ (.D(_0120_),
    .RN(net34),
    .CLK(clknet_leaf_47_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4959_ (.D(_0121_),
    .RN(net34),
    .CLK(clknet_leaf_46_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4960_ (.D(_0122_),
    .RN(net34),
    .CLK(clknet_leaf_47_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4961_ (.D(_0123_),
    .RN(net34),
    .CLK(clknet_leaf_30_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4962_ (.D(_0124_),
    .RN(net34),
    .CLK(clknet_leaf_30_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4963_ (.D(_0125_),
    .RN(net34),
    .CLK(clknet_leaf_31_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4964_ (.D(_0126_),
    .RN(net34),
    .CLK(clknet_leaf_30_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4965_ (.D(_0127_),
    .RN(net34),
    .CLK(clknet_leaf_38_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4966_ (.D(_0128_),
    .RN(net34),
    .CLK(clknet_leaf_38_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4967_ (.D(_0129_),
    .RN(net34),
    .CLK(clknet_leaf_38_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4968_ (.D(_0130_),
    .RN(net34),
    .CLK(clknet_leaf_38_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4969_ (.D(_0131_),
    .RN(net34),
    .CLK(clknet_leaf_40_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4970_ (.D(_0132_),
    .RN(net34),
    .CLK(clknet_leaf_41_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4971_ (.D(_0133_),
    .RN(net34),
    .CLK(clknet_leaf_41_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4972_ (.D(_0134_),
    .RN(net34),
    .CLK(clknet_leaf_50_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4973_ (.D(_0135_),
    .RN(net34),
    .CLK(clknet_leaf_46_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4974_ (.D(_0136_),
    .RN(net34),
    .CLK(clknet_leaf_47_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4975_ (.D(_0137_),
    .RN(net34),
    .CLK(clknet_leaf_47_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4976_ (.D(_0138_),
    .RN(net34),
    .CLK(clknet_leaf_46_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4977_ (.D(_0139_),
    .RN(net34),
    .CLK(clknet_leaf_25_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4978_ (.D(_0140_),
    .RN(net34),
    .CLK(clknet_leaf_23_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4979_ (.D(_0141_),
    .RN(net34),
    .CLK(clknet_leaf_23_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4980_ (.D(_0142_),
    .RN(net34),
    .CLK(clknet_leaf_24_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4981_ (.D(_0143_),
    .RN(net34),
    .CLK(clknet_leaf_63_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4982_ (.D(_0144_),
    .RN(net34),
    .CLK(clknet_leaf_63_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4983_ (.D(_0145_),
    .RN(net34),
    .CLK(clknet_leaf_63_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4984_ (.D(_0146_),
    .RN(net34),
    .CLK(clknet_leaf_63_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4985_ (.D(_0147_),
    .RN(net34),
    .CLK(clknet_leaf_60_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4986_ (.D(_0148_),
    .RN(net34),
    .CLK(clknet_leaf_60_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4987_ (.D(_0149_),
    .RN(net34),
    .CLK(clknet_leaf_51_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4988_ (.D(_0150_),
    .RN(net34),
    .CLK(clknet_leaf_60_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4989_ (.D(_0151_),
    .RN(net34),
    .CLK(clknet_leaf_56_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4990_ (.D(_0152_),
    .RN(net34),
    .CLK(clknet_leaf_55_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4991_ (.D(_0153_),
    .RN(net34),
    .CLK(clknet_leaf_55_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4992_ (.D(_0154_),
    .RN(net34),
    .CLK(clknet_leaf_55_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4993_ (.D(_0155_),
    .RN(net34),
    .CLK(clknet_leaf_23_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4994_ (.D(_0156_),
    .RN(net34),
    .CLK(clknet_leaf_23_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4995_ (.D(_0157_),
    .RN(net34),
    .CLK(clknet_leaf_23_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4996_ (.D(_0158_),
    .RN(net34),
    .CLK(clknet_leaf_23_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4997_ (.D(_0159_),
    .RN(net34),
    .CLK(clknet_leaf_65_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4998_ (.D(_0160_),
    .RN(net34),
    .CLK(clknet_leaf_65_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _4999_ (.D(_0161_),
    .RN(net34),
    .CLK(clknet_leaf_65_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5000_ (.D(_0162_),
    .RN(net34),
    .CLK(clknet_leaf_64_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5001_ (.D(_0163_),
    .RN(net34),
    .CLK(clknet_leaf_57_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5002_ (.D(_0164_),
    .RN(net34),
    .CLK(clknet_leaf_57_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5003_ (.D(_0165_),
    .RN(net34),
    .CLK(clknet_leaf_57_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5004_ (.D(_0166_),
    .RN(net34),
    .CLK(clknet_leaf_59_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5005_ (.D(_0167_),
    .RN(net34),
    .CLK(clknet_leaf_55_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5006_ (.D(_0168_),
    .RN(net34),
    .CLK(clknet_leaf_55_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5007_ (.D(_0169_),
    .RN(net34),
    .CLK(clknet_leaf_55_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5008_ (.D(_0170_),
    .RN(net34),
    .CLK(clknet_leaf_55_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5009_ (.D(_0171_),
    .RN(net34),
    .CLK(clknet_leaf_121_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5010_ (.D(_0172_),
    .RN(net34),
    .CLK(clknet_leaf_109_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5011_ (.D(_0173_),
    .RN(net34),
    .CLK(clknet_leaf_121_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5012_ (.D(_0174_),
    .RN(net34),
    .CLK(clknet_leaf_67_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5013_ (.D(_0175_),
    .RN(net34),
    .CLK(clknet_leaf_68_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5014_ (.D(_0176_),
    .RN(net34),
    .CLK(clknet_leaf_68_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5015_ (.D(_0177_),
    .RN(net34),
    .CLK(clknet_leaf_69_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5016_ (.D(_0178_),
    .RN(net34),
    .CLK(clknet_leaf_69_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5017_ (.D(_0179_),
    .RN(net34),
    .CLK(clknet_leaf_58_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5018_ (.D(_0180_),
    .RN(net34),
    .CLK(clknet_leaf_58_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5019_ (.D(_0181_),
    .RN(net34),
    .CLK(clknet_leaf_58_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5020_ (.D(_0182_),
    .RN(net34),
    .CLK(clknet_leaf_75_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5021_ (.D(_0183_),
    .RN(net34),
    .CLK(clknet_leaf_77_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5022_ (.D(_0184_),
    .RN(net34),
    .CLK(clknet_leaf_55_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5023_ (.D(_0185_),
    .RN(net34),
    .CLK(clknet_leaf_77_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5024_ (.D(_0186_),
    .RN(net34),
    .CLK(clknet_leaf_55_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5025_ (.D(_0187_),
    .RN(net34),
    .CLK(clknet_leaf_108_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5026_ (.D(_0188_),
    .RN(net34),
    .CLK(clknet_leaf_109_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5027_ (.D(_0189_),
    .RN(net34),
    .CLK(clknet_leaf_109_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5028_ (.D(_0190_),
    .RN(net34),
    .CLK(clknet_leaf_108_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5029_ (.D(_0191_),
    .RN(net34),
    .CLK(clknet_leaf_68_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5030_ (.D(_0192_),
    .RN(net34),
    .CLK(clknet_leaf_69_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5031_ (.D(_0193_),
    .RN(net34),
    .CLK(clknet_leaf_69_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5032_ (.D(_0194_),
    .RN(net34),
    .CLK(clknet_leaf_65_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5033_ (.D(_0195_),
    .RN(net34),
    .CLK(clknet_leaf_57_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5034_ (.D(_0196_),
    .RN(net34),
    .CLK(clknet_leaf_75_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5035_ (.D(_0197_),
    .RN(net34),
    .CLK(clknet_leaf_58_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5036_ (.D(_0198_),
    .RN(net34),
    .CLK(clknet_leaf_58_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5037_ (.D(_0199_),
    .RN(net34),
    .CLK(clknet_leaf_77_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5038_ (.D(_0200_),
    .RN(net34),
    .CLK(clknet_leaf_77_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5039_ (.D(_0201_),
    .RN(net34),
    .CLK(clknet_leaf_77_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5040_ (.D(_0202_),
    .RN(net34),
    .CLK(clknet_leaf_77_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5041_ (.D(_0203_),
    .RN(net34),
    .CLK(clknet_leaf_106_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5042_ (.D(_0204_),
    .RN(net34),
    .CLK(clknet_leaf_105_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5043_ (.D(_0205_),
    .RN(net34),
    .CLK(clknet_4_0_0_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5044_ (.D(_0206_),
    .RN(net34),
    .CLK(clknet_leaf_105_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5045_ (.D(_0207_),
    .RN(net34),
    .CLK(clknet_leaf_103_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5046_ (.D(_0208_),
    .RN(net34),
    .CLK(clknet_leaf_103_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5047_ (.D(_0209_),
    .RN(net34),
    .CLK(clknet_leaf_103_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5048_ (.D(_0210_),
    .RN(net34),
    .CLK(clknet_leaf_103_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5049_ (.D(_0211_),
    .RN(net34),
    .CLK(clknet_leaf_73_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5050_ (.D(_0212_),
    .RN(net34),
    .CLK(clknet_leaf_102_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5051_ (.D(_0213_),
    .RN(net34),
    .CLK(clknet_leaf_91_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5052_ (.D(_0214_),
    .RN(net34),
    .CLK(clknet_leaf_73_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5053_ (.D(_0215_),
    .RN(net34),
    .CLK(clknet_leaf_78_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5054_ (.D(_0216_),
    .RN(net34),
    .CLK(clknet_leaf_78_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5055_ (.D(_0217_),
    .RN(net34),
    .CLK(clknet_leaf_78_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5056_ (.D(_0218_),
    .RN(net34),
    .CLK(clknet_leaf_79_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5057_ (.D(_0219_),
    .RN(net34),
    .CLK(clknet_leaf_99_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5058_ (.D(_0220_),
    .RN(net34),
    .CLK(clknet_leaf_99_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5059_ (.D(_0221_),
    .RN(net34),
    .CLK(clknet_leaf_100_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5060_ (.D(_0222_),
    .RN(net34),
    .CLK(clknet_leaf_100_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5061_ (.D(_0223_),
    .RN(net34),
    .CLK(clknet_leaf_100_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5062_ (.D(_0224_),
    .RN(net34),
    .CLK(clknet_leaf_100_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5063_ (.D(_0225_),
    .RN(net34),
    .CLK(clknet_leaf_101_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5064_ (.D(_0226_),
    .RN(net34),
    .CLK(clknet_leaf_101_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5065_ (.D(_0227_),
    .RN(net34),
    .CLK(clknet_leaf_73_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5066_ (.D(_0228_),
    .RN(net34),
    .CLK(clknet_leaf_91_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5067_ (.D(_0229_),
    .RN(net34),
    .CLK(clknet_leaf_83_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5068_ (.D(_0230_),
    .RN(net34),
    .CLK(clknet_leaf_91_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5069_ (.D(_0231_),
    .RN(net34),
    .CLK(clknet_leaf_81_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5070_ (.D(_0232_),
    .RN(net34),
    .CLK(clknet_leaf_80_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5071_ (.D(_0233_),
    .RN(net34),
    .CLK(clknet_leaf_80_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5072_ (.D(_0234_),
    .RN(net34),
    .CLK(clknet_leaf_80_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5073_ (.D(_0235_),
    .RN(net34),
    .CLK(clknet_leaf_105_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5074_ (.D(_0236_),
    .RN(net34),
    .CLK(clknet_leaf_105_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5075_ (.D(_0237_),
    .RN(net34),
    .CLK(clknet_leaf_105_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5076_ (.D(_0238_),
    .RN(net34),
    .CLK(clknet_leaf_104_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5077_ (.D(_0239_),
    .RN(net34),
    .CLK(clknet_leaf_104_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5078_ (.D(_0240_),
    .RN(net34),
    .CLK(clknet_leaf_104_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5079_ (.D(_0241_),
    .RN(net34),
    .CLK(clknet_leaf_103_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5080_ (.D(_0242_),
    .RN(net34),
    .CLK(clknet_leaf_102_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5081_ (.D(_0243_),
    .RN(net34),
    .CLK(clknet_leaf_73_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5082_ (.D(_0244_),
    .RN(net34),
    .CLK(clknet_leaf_82_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5083_ (.D(_0245_),
    .RN(net34),
    .CLK(clknet_leaf_83_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5084_ (.D(_0246_),
    .RN(net34),
    .CLK(clknet_leaf_83_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5085_ (.D(_0247_),
    .RN(net34),
    .CLK(clknet_leaf_79_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5086_ (.D(_0248_),
    .RN(net34),
    .CLK(clknet_leaf_78_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5087_ (.D(_0249_),
    .RN(net34),
    .CLK(clknet_leaf_78_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5088_ (.D(_0250_),
    .RN(net34),
    .CLK(clknet_leaf_78_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5089_ (.D(_0251_),
    .RN(net34),
    .CLK(clknet_leaf_115_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5090_ (.D(_0252_),
    .RN(net34),
    .CLK(clknet_leaf_116_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5091_ (.D(_0253_),
    .RN(net34),
    .CLK(clknet_leaf_99_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5092_ (.D(_0254_),
    .RN(net34),
    .CLK(clknet_leaf_100_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5093_ (.D(_0255_),
    .RN(net34),
    .CLK(clknet_leaf_100_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5094_ (.D(_0256_),
    .RN(net34),
    .CLK(clknet_leaf_100_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5095_ (.D(_0257_),
    .RN(net34),
    .CLK(clknet_leaf_102_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5096_ (.D(_0258_),
    .RN(net34),
    .CLK(clknet_leaf_101_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5097_ (.D(_0259_),
    .RN(net34),
    .CLK(clknet_leaf_82_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5098_ (.D(_0260_),
    .RN(net34),
    .CLK(clknet_leaf_91_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5099_ (.D(_0261_),
    .RN(net34),
    .CLK(clknet_leaf_91_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5100_ (.D(_0262_),
    .RN(net34),
    .CLK(clknet_leaf_91_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5101_ (.D(_0263_),
    .RN(net34),
    .CLK(clknet_leaf_81_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5102_ (.D(_0264_),
    .RN(net34),
    .CLK(clknet_leaf_80_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5103_ (.D(_0265_),
    .RN(net34),
    .CLK(clknet_leaf_79_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5104_ (.D(_0266_),
    .RN(net34),
    .CLK(clknet_leaf_80_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5105_ (.D(_0267_),
    .RN(net34),
    .CLK(clknet_leaf_115_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5106_ (.D(_0268_),
    .RN(net34),
    .CLK(clknet_leaf_115_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5107_ (.D(_0269_),
    .RN(net34),
    .CLK(clknet_leaf_115_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5108_ (.D(_0270_),
    .RN(net34),
    .CLK(clknet_leaf_115_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5109_ (.D(_0271_),
    .RN(net34),
    .CLK(clknet_leaf_101_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5110_ (.D(_0272_),
    .RN(net34),
    .CLK(clknet_leaf_96_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5111_ (.D(_0273_),
    .RN(net34),
    .CLK(clknet_leaf_94_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5112_ (.D(_0274_),
    .RN(net34),
    .CLK(clknet_leaf_94_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5113_ (.D(_0275_),
    .RN(net34),
    .CLK(clknet_leaf_90_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5114_ (.D(_0276_),
    .RN(net34),
    .CLK(clknet_leaf_87_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5115_ (.D(_0277_),
    .RN(net34),
    .CLK(clknet_leaf_83_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5116_ (.D(_0278_),
    .RN(net34),
    .CLK(clknet_leaf_90_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5117_ (.D(_0279_),
    .RN(net34),
    .CLK(clknet_leaf_84_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5118_ (.D(_0280_),
    .RN(net34),
    .CLK(clknet_leaf_86_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5119_ (.D(_0281_),
    .RN(net34),
    .CLK(clknet_leaf_85_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5120_ (.D(_0282_),
    .RN(net34),
    .CLK(clknet_leaf_85_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5121_ (.D(_0283_),
    .RN(net34),
    .CLK(clknet_leaf_117_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5122_ (.D(_0284_),
    .RN(net34),
    .CLK(clknet_leaf_116_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5123_ (.D(_0285_),
    .RN(net34),
    .CLK(clknet_leaf_116_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5124_ (.D(_0286_),
    .RN(net34),
    .CLK(clknet_leaf_117_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5125_ (.D(_0287_),
    .RN(net34),
    .CLK(clknet_leaf_101_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5126_ (.D(_0288_),
    .RN(net34),
    .CLK(clknet_leaf_94_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5127_ (.D(_0289_),
    .RN(net34),
    .CLK(clknet_leaf_94_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5128_ (.D(_0290_),
    .RN(net34),
    .CLK(clknet_leaf_92_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5129_ (.D(_0291_),
    .RN(net34),
    .CLK(clknet_leaf_87_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5130_ (.D(_0292_),
    .RN(net34),
    .CLK(clknet_leaf_88_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5131_ (.D(_0293_),
    .RN(net34),
    .CLK(clknet_leaf_90_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5132_ (.D(_0294_),
    .RN(net34),
    .CLK(clknet_leaf_88_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5133_ (.D(_0295_),
    .RN(net34),
    .CLK(clknet_leaf_86_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5134_ (.D(_0296_),
    .RN(net34),
    .CLK(clknet_leaf_86_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5135_ (.D(_0297_),
    .RN(net34),
    .CLK(clknet_leaf_85_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5136_ (.D(_0298_),
    .RN(net34),
    .CLK(clknet_leaf_85_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5137_ (.D(_0299_),
    .RN(net34),
    .CLK(clknet_leaf_117_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5138_ (.D(_0300_),
    .RN(net34),
    .CLK(clknet_leaf_114_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5139_ (.D(_0301_),
    .RN(net34),
    .CLK(clknet_leaf_114_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5140_ (.D(_0302_),
    .RN(net34),
    .CLK(clknet_leaf_117_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5141_ (.D(_0303_),
    .RN(net34),
    .CLK(clknet_leaf_101_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5142_ (.D(_0304_),
    .RN(net34),
    .CLK(clknet_leaf_96_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5143_ (.D(_0305_),
    .RN(net34),
    .CLK(clknet_leaf_94_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5144_ (.D(_0306_),
    .RN(net34),
    .CLK(clknet_leaf_94_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5145_ (.D(_0307_),
    .RN(net34),
    .CLK(clknet_leaf_87_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5146_ (.D(_0308_),
    .RN(net34),
    .CLK(clknet_leaf_87_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5147_ (.D(_0309_),
    .RN(net34),
    .CLK(clknet_leaf_90_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5148_ (.D(_0310_),
    .RN(net34),
    .CLK(clknet_leaf_87_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5149_ (.D(_0311_),
    .RN(net34),
    .CLK(clknet_leaf_84_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5150_ (.D(_0312_),
    .RN(net34),
    .CLK(clknet_leaf_86_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5151_ (.D(_0313_),
    .RN(net34),
    .CLK(clknet_leaf_85_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5152_ (.D(_0314_),
    .RN(net34),
    .CLK(clknet_leaf_85_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5153_ (.D(_0315_),
    .RN(net34),
    .CLK(clknet_leaf_117_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5154_ (.D(_0316_),
    .RN(net34),
    .CLK(clknet_leaf_114_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5155_ (.D(_0317_),
    .RN(net34),
    .CLK(clknet_leaf_114_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5156_ (.D(_0318_),
    .RN(net34),
    .CLK(clknet_leaf_116_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5157_ (.D(_0319_),
    .RN(net34),
    .CLK(clknet_leaf_101_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5158_ (.D(_0320_),
    .RN(net34),
    .CLK(clknet_leaf_94_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5159_ (.D(_0321_),
    .RN(net34),
    .CLK(clknet_leaf_94_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5160_ (.D(_0322_),
    .RN(net34),
    .CLK(clknet_leaf_92_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5161_ (.D(_0323_),
    .RN(net34),
    .CLK(clknet_leaf_87_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5162_ (.D(_0324_),
    .RN(net34),
    .CLK(clknet_leaf_87_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5163_ (.D(_0325_),
    .RN(net34),
    .CLK(clknet_leaf_90_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5164_ (.D(_0326_),
    .RN(net34),
    .CLK(clknet_leaf_87_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5165_ (.D(_0327_),
    .RN(net34),
    .CLK(clknet_leaf_86_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5166_ (.D(_0328_),
    .RN(net34),
    .CLK(clknet_leaf_86_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5167_ (.D(_0329_),
    .RN(net34),
    .CLK(clknet_leaf_85_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5168_ (.D(_0330_),
    .RN(net34),
    .CLK(clknet_leaf_85_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5169_ (.D(_0331_),
    .RN(net34),
    .CLK(clknet_leaf_114_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5170_ (.D(_0332_),
    .RN(net34),
    .CLK(clknet_leaf_114_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5171_ (.D(_0333_),
    .RN(net34),
    .CLK(clknet_leaf_114_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5172_ (.D(_0334_),
    .RN(net34),
    .CLK(clknet_leaf_112_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5173_ (.D(_0335_),
    .RN(net34),
    .CLK(clknet_leaf_98_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5174_ (.D(_0336_),
    .RN(net34),
    .CLK(clknet_4_8_0_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5175_ (.D(_0337_),
    .RN(net34),
    .CLK(clknet_leaf_96_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5176_ (.D(_0338_),
    .RN(net34),
    .CLK(clknet_leaf_98_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5177_ (.D(_0339_),
    .RN(net34),
    .CLK(clknet_leaf_93_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5178_ (.D(_0340_),
    .RN(net34),
    .CLK(clknet_leaf_93_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5179_ (.D(_0341_),
    .RN(net34),
    .CLK(clknet_4_10_0_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5180_ (.D(_0342_),
    .RN(net34),
    .CLK(clknet_leaf_88_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5181_ (.D(_0343_),
    .RN(net34),
    .CLK(clknet_leaf_72_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5182_ (.D(_0344_),
    .RN(net34),
    .CLK(clknet_leaf_81_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5183_ (.D(_0345_),
    .RN(net34),
    .CLK(clknet_leaf_84_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5184_ (.D(_0346_),
    .RN(net34),
    .CLK(clknet_leaf_83_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5185_ (.D(_0347_),
    .RN(net34),
    .CLK(clknet_leaf_112_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5186_ (.D(_0348_),
    .RN(net34),
    .CLK(clknet_leaf_112_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5187_ (.D(_0349_),
    .RN(net34),
    .CLK(clknet_leaf_113_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5188_ (.D(_0350_),
    .RN(net34),
    .CLK(clknet_leaf_112_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5189_ (.D(_0351_),
    .RN(net34),
    .CLK(clknet_leaf_98_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5190_ (.D(_0352_),
    .RN(net34),
    .CLK(clknet_leaf_96_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5191_ (.D(_0353_),
    .RN(net34),
    .CLK(clknet_leaf_96_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5192_ (.D(_0354_),
    .RN(net34),
    .CLK(clknet_leaf_97_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5193_ (.D(_0355_),
    .RN(net34),
    .CLK(clknet_leaf_92_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5194_ (.D(_0356_),
    .RN(net34),
    .CLK(clknet_leaf_93_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5195_ (.D(_0357_),
    .RN(net34),
    .CLK(clknet_leaf_92_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5196_ (.D(_0358_),
    .RN(net34),
    .CLK(clknet_leaf_92_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5197_ (.D(_0359_),
    .RN(net34),
    .CLK(clknet_leaf_102_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5198_ (.D(_0360_),
    .RN(net34),
    .CLK(clknet_leaf_82_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5199_ (.D(_0361_),
    .RN(net34),
    .CLK(clknet_leaf_81_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5200_ (.D(_0362_),
    .RN(net34),
    .CLK(clknet_leaf_84_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5201_ (.D(_0363_),
    .RN(net34),
    .CLK(clknet_leaf_113_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5202_ (.D(_0364_),
    .RN(net34),
    .CLK(clknet_leaf_113_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5203_ (.D(_0365_),
    .RN(net34),
    .CLK(clknet_leaf_113_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5204_ (.D(_0366_),
    .RN(net34),
    .CLK(clknet_leaf_110_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5205_ (.D(_0367_),
    .RN(net34),
    .CLK(clknet_leaf_98_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5206_ (.D(_0368_),
    .RN(net34),
    .CLK(clknet_leaf_97_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5207_ (.D(_0369_),
    .RN(net34),
    .CLK(clknet_leaf_96_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5208_ (.D(_0370_),
    .RN(net34),
    .CLK(clknet_leaf_97_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5209_ (.D(_0371_),
    .RN(net34),
    .CLK(clknet_leaf_92_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5210_ (.D(_0372_),
    .RN(net34),
    .CLK(clknet_leaf_93_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5211_ (.D(_0373_),
    .RN(net34),
    .CLK(clknet_leaf_91_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5212_ (.D(_0374_),
    .RN(net34),
    .CLK(clknet_leaf_102_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5213_ (.D(_0375_),
    .RN(net34),
    .CLK(clknet_leaf_72_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5214_ (.D(_0376_),
    .RN(net34),
    .CLK(clknet_leaf_82_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5215_ (.D(_0377_),
    .RN(net34),
    .CLK(clknet_leaf_81_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5216_ (.D(_0378_),
    .RN(net34),
    .CLK(clknet_leaf_84_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5217_ (.D(_0379_),
    .RN(net34),
    .CLK(clknet_leaf_113_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5218_ (.D(_0380_),
    .RN(net34),
    .CLK(clknet_leaf_113_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5219_ (.D(_0381_),
    .RN(net34),
    .CLK(clknet_leaf_113_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5220_ (.D(_0382_),
    .RN(net34),
    .CLK(clknet_leaf_110_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5221_ (.D(_0383_),
    .RN(net34),
    .CLK(clknet_leaf_98_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5222_ (.D(_0384_),
    .RN(net34),
    .CLK(clknet_leaf_97_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5223_ (.D(_0385_),
    .RN(net34),
    .CLK(clknet_leaf_96_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5224_ (.D(_0386_),
    .RN(net34),
    .CLK(clknet_leaf_97_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5225_ (.D(_0387_),
    .RN(net34),
    .CLK(clknet_leaf_93_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5226_ (.D(_0388_),
    .RN(net34),
    .CLK(clknet_leaf_93_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5227_ (.D(_0389_),
    .RN(net34),
    .CLK(clknet_leaf_91_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5228_ (.D(_0390_),
    .RN(net34),
    .CLK(clknet_leaf_91_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5229_ (.D(_0391_),
    .RN(net34),
    .CLK(clknet_leaf_72_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5230_ (.D(_0392_),
    .RN(net34),
    .CLK(clknet_leaf_82_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5231_ (.D(_0393_),
    .RN(net34),
    .CLK(clknet_leaf_81_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5232_ (.D(_0394_),
    .RN(net34),
    .CLK(clknet_leaf_84_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5233_ (.D(_0395_),
    .RN(net34),
    .CLK(clknet_leaf_110_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5234_ (.D(_0396_),
    .RN(net34),
    .CLK(clknet_leaf_118_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5235_ (.D(_0397_),
    .RN(net34),
    .CLK(clknet_leaf_118_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5236_ (.D(_0398_),
    .RN(net34),
    .CLK(clknet_leaf_110_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5237_ (.D(_0399_),
    .RN(net34),
    .CLK(clknet_leaf_106_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5238_ (.D(_0400_),
    .RN(net34),
    .CLK(clknet_leaf_106_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5239_ (.D(_0401_),
    .RN(net34),
    .CLK(clknet_leaf_104_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5240_ (.D(_0402_),
    .RN(net34),
    .CLK(clknet_leaf_106_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5241_ (.D(_0403_),
    .RN(net34),
    .CLK(clknet_leaf_72_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5242_ (.D(_0404_),
    .RN(net34),
    .CLK(clknet_leaf_71_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5243_ (.D(_0405_),
    .RN(net34),
    .CLK(clknet_leaf_72_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5244_ (.D(_0406_),
    .RN(net34),
    .CLK(clknet_leaf_72_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5245_ (.D(_0407_),
    .RN(net34),
    .CLK(clknet_leaf_73_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5246_ (.D(_0408_),
    .RN(net34),
    .CLK(clknet_leaf_73_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5247_ (.D(_0409_),
    .RN(net34),
    .CLK(clknet_leaf_74_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5248_ (.D(_0410_),
    .RN(net34),
    .CLK(clknet_leaf_74_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5249_ (.D(_0411_),
    .RN(net34),
    .CLK(clknet_leaf_120_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5250_ (.D(_0412_),
    .RN(net34),
    .CLK(clknet_leaf_119_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5251_ (.D(_0413_),
    .RN(net34),
    .CLK(clknet_leaf_119_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5252_ (.D(_0414_),
    .RN(net34),
    .CLK(clknet_leaf_110_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5253_ (.D(_0415_),
    .RN(net34),
    .CLK(clknet_leaf_67_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5254_ (.D(_0416_),
    .RN(net34),
    .CLK(clknet_leaf_106_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5255_ (.D(_0417_),
    .RN(net34),
    .CLK(clknet_leaf_68_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5256_ (.D(_0418_),
    .RN(net34),
    .CLK(clknet_leaf_71_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5257_ (.D(_0419_),
    .RN(net34),
    .CLK(clknet_leaf_70_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5258_ (.D(_0420_),
    .RN(net34),
    .CLK(clknet_leaf_71_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5259_ (.D(_0421_),
    .RN(net34),
    .CLK(clknet_leaf_70_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5260_ (.D(_0422_),
    .RN(net34),
    .CLK(clknet_leaf_70_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5261_ (.D(_0423_),
    .RN(net34),
    .CLK(clknet_leaf_74_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5262_ (.D(_0424_),
    .RN(net34),
    .CLK(clknet_leaf_74_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5263_ (.D(_0425_),
    .RN(net34),
    .CLK(clknet_leaf_76_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5264_ (.D(_0426_),
    .RN(net34),
    .CLK(clknet_leaf_78_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5265_ (.D(_0427_),
    .RN(net34),
    .CLK(clknet_leaf_120_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5266_ (.D(_0428_),
    .RN(net34),
    .CLK(clknet_leaf_120_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5267_ (.D(_0429_),
    .RN(net34),
    .CLK(clknet_leaf_118_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5268_ (.D(_0430_),
    .RN(net34),
    .CLK(clknet_leaf_120_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5269_ (.D(_0431_),
    .RN(net34),
    .CLK(clknet_leaf_108_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5270_ (.D(_0432_),
    .RN(net34),
    .CLK(clknet_leaf_107_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5271_ (.D(_0433_),
    .RN(net34),
    .CLK(clknet_leaf_68_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5272_ (.D(_0434_),
    .RN(net34),
    .CLK(clknet_leaf_107_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5273_ (.D(_0435_),
    .RN(net34),
    .CLK(clknet_leaf_70_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5274_ (.D(_0436_),
    .RN(net34),
    .CLK(clknet_leaf_71_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5275_ (.D(_0437_),
    .RN(net34),
    .CLK(clknet_leaf_70_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5276_ (.D(_0438_),
    .RN(net34),
    .CLK(clknet_leaf_69_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5277_ (.D(_0439_),
    .RN(net34),
    .CLK(clknet_leaf_75_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5278_ (.D(_0440_),
    .RN(net34),
    .CLK(clknet_leaf_76_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5279_ (.D(_0441_),
    .RN(net34),
    .CLK(clknet_leaf_76_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5280_ (.D(_0442_),
    .RN(net34),
    .CLK(clknet_leaf_76_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5281_ (.D(_0443_),
    .RN(net34),
    .CLK(clknet_leaf_120_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5282_ (.D(_0444_),
    .RN(net34),
    .CLK(clknet_leaf_119_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5283_ (.D(_0445_),
    .RN(net34),
    .CLK(clknet_leaf_118_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5284_ (.D(_0446_),
    .RN(net34),
    .CLK(clknet_leaf_109_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5285_ (.D(_0447_),
    .RN(net34),
    .CLK(clknet_leaf_67_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5286_ (.D(_0448_),
    .RN(net34),
    .CLK(clknet_leaf_107_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5287_ (.D(_0449_),
    .RN(net34),
    .CLK(clknet_leaf_68_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5288_ (.D(_0450_),
    .RN(net34),
    .CLK(clknet_leaf_68_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5289_ (.D(_0451_),
    .RN(net34),
    .CLK(clknet_leaf_70_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5290_ (.D(_0452_),
    .RN(net34),
    .CLK(clknet_leaf_71_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5291_ (.D(_0453_),
    .RN(net34),
    .CLK(clknet_leaf_70_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5292_ (.D(_0454_),
    .RN(net34),
    .CLK(clknet_leaf_69_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5293_ (.D(_0455_),
    .RN(net34),
    .CLK(clknet_leaf_75_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5294_ (.D(_0456_),
    .RN(net34),
    .CLK(clknet_leaf_76_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5295_ (.D(_0457_),
    .RN(net34),
    .CLK(clknet_leaf_76_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5296_ (.D(_0458_),
    .RN(net34),
    .CLK(clknet_leaf_76_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5297_ (.D(_0459_),
    .RN(net34),
    .CLK(clknet_leaf_0_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5298_ (.D(_0460_),
    .RN(net34),
    .CLK(clknet_leaf_2_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5299_ (.D(_0461_),
    .RN(net34),
    .CLK(clknet_leaf_2_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5300_ (.D(_0462_),
    .RN(net34),
    .CLK(clknet_leaf_121_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5301_ (.D(_0463_),
    .RN(net34),
    .CLK(clknet_leaf_67_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5302_ (.D(_0464_),
    .RN(net34),
    .CLK(clknet_leaf_67_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5303_ (.D(_0465_),
    .RN(net34),
    .CLK(clknet_leaf_67_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5304_ (.D(_0466_),
    .RN(net34),
    .CLK(clknet_leaf_67_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5305_ (.D(_0467_),
    .RN(net34),
    .CLK(clknet_leaf_64_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5306_ (.D(_0468_),
    .RN(net34),
    .CLK(clknet_leaf_64_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5307_ (.D(_0469_),
    .RN(net34),
    .CLK(clknet_leaf_64_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5308_ (.D(_0470_),
    .RN(net34),
    .CLK(clknet_leaf_64_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5309_ (.D(_0471_),
    .RN(net34),
    .CLK(clknet_leaf_57_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5310_ (.D(_0472_),
    .RN(net34),
    .CLK(clknet_leaf_56_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5311_ (.D(_0473_),
    .RN(net34),
    .CLK(clknet_leaf_54_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5312_ (.D(_0474_),
    .RN(net34),
    .CLK(clknet_leaf_54_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5313_ (.D(_0475_),
    .RN(net34),
    .CLK(clknet_leaf_0_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5314_ (.D(_0476_),
    .RN(net34),
    .CLK(clknet_leaf_1_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5315_ (.D(_0477_),
    .RN(net34),
    .CLK(clknet_leaf_1_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5316_ (.D(_0478_),
    .RN(net34),
    .CLK(clknet_leaf_0_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5317_ (.D(_0479_),
    .RN(net34),
    .CLK(clknet_leaf_66_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5318_ (.D(_0480_),
    .RN(net34),
    .CLK(clknet_leaf_24_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5319_ (.D(_0481_),
    .RN(net34),
    .CLK(clknet_leaf_66_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5320_ (.D(_0482_),
    .RN(net34),
    .CLK(clknet_leaf_66_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5321_ (.D(_0483_),
    .RN(net34),
    .CLK(clknet_leaf_59_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5322_ (.D(_0484_),
    .RN(net34),
    .CLK(clknet_leaf_64_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5323_ (.D(_0485_),
    .RN(net34),
    .CLK(clknet_leaf_59_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5324_ (.D(_0486_),
    .RN(net34),
    .CLK(clknet_leaf_59_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5325_ (.D(_0487_),
    .RN(net34),
    .CLK(clknet_leaf_57_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5326_ (.D(_0488_),
    .RN(net34),
    .CLK(clknet_leaf_54_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5327_ (.D(_0489_),
    .RN(net34),
    .CLK(clknet_leaf_54_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5328_ (.D(_0490_),
    .RN(net34),
    .CLK(clknet_leaf_54_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5329_ (.D(_0491_),
    .RN(net34),
    .CLK(clknet_leaf_0_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5330_ (.D(_0492_),
    .RN(net34),
    .CLK(clknet_leaf_1_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5331_ (.D(_0493_),
    .RN(net34),
    .CLK(clknet_leaf_0_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5332_ (.D(_0494_),
    .RN(net34),
    .CLK(clknet_leaf_0_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5333_ (.D(_0495_),
    .RN(net34),
    .CLK(clknet_leaf_66_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5334_ (.D(_0496_),
    .RN(net34),
    .CLK(clknet_leaf_23_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5335_ (.D(_0497_),
    .RN(net34),
    .CLK(clknet_leaf_66_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5336_ (.D(_0498_),
    .RN(net34),
    .CLK(clknet_leaf_66_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5337_ (.D(_0499_),
    .RN(net34),
    .CLK(clknet_leaf_59_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5338_ (.D(_0500_),
    .RN(net34),
    .CLK(clknet_leaf_62_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5339_ (.D(_0501_),
    .RN(net34),
    .CLK(clknet_leaf_59_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5340_ (.D(_0502_),
    .RN(net34),
    .CLK(clknet_leaf_60_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5341_ (.D(_0503_),
    .RN(net34),
    .CLK(clknet_leaf_51_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5342_ (.D(_0504_),
    .RN(net34),
    .CLK(clknet_leaf_53_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5343_ (.D(_0505_),
    .RN(net34),
    .CLK(clknet_leaf_54_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5344_ (.D(_0506_),
    .RN(net34),
    .CLK(clknet_leaf_53_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5345_ (.D(_0507_),
    .RN(net34),
    .CLK(clknet_leaf_1_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5346_ (.D(_0508_),
    .RN(net34),
    .CLK(clknet_leaf_3_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5347_ (.D(_0509_),
    .RN(net34),
    .CLK(clknet_leaf_3_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5348_ (.D(_0510_),
    .RN(net34),
    .CLK(clknet_leaf_22_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5349_ (.D(_0511_),
    .RN(net34),
    .CLK(clknet_leaf_27_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5350_ (.D(_0512_),
    .RN(net34),
    .CLK(clknet_leaf_24_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5351_ (.D(_0513_),
    .RN(net34),
    .CLK(clknet_leaf_24_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5352_ (.D(_0514_),
    .RN(net34),
    .CLK(clknet_leaf_24_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5353_ (.D(_0515_),
    .RN(net34),
    .CLK(clknet_leaf_61_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5354_ (.D(_0516_),
    .RN(net34),
    .CLK(clknet_leaf_61_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5355_ (.D(_0517_),
    .RN(net34),
    .CLK(clknet_leaf_61_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5356_ (.D(_0518_),
    .RN(net34),
    .CLK(clknet_leaf_60_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5357_ (.D(_0519_),
    .RN(net34),
    .CLK(clknet_leaf_51_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5358_ (.D(_0520_),
    .RN(net34),
    .CLK(clknet_leaf_52_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5359_ (.D(_0521_),
    .RN(net34),
    .CLK(clknet_leaf_53_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5360_ (.D(_0522_),
    .RN(net34),
    .CLK(clknet_leaf_52_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5361_ (.D(_0523_),
    .RN(net34),
    .CLK(clknet_leaf_22_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5362_ (.D(_0524_),
    .RN(net34),
    .CLK(clknet_leaf_22_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5363_ (.D(_0525_),
    .RN(net34),
    .CLK(clknet_leaf_22_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5364_ (.D(_0526_),
    .RN(net34),
    .CLK(clknet_leaf_22_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5365_ (.D(_0527_),
    .RN(net34),
    .CLK(clknet_leaf_27_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5366_ (.D(_0528_),
    .RN(net34),
    .CLK(clknet_leaf_27_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5367_ (.D(_0529_),
    .RN(net34),
    .CLK(clknet_leaf_62_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5368_ (.D(_0530_),
    .RN(net34),
    .CLK(clknet_leaf_62_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5369_ (.D(_0531_),
    .RN(net34),
    .CLK(clknet_leaf_51_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5370_ (.D(_0532_),
    .RN(net34),
    .CLK(clknet_leaf_51_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5371_ (.D(_0533_),
    .RN(net34),
    .CLK(clknet_leaf_61_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5372_ (.D(_0534_),
    .RN(net34),
    .CLK(clknet_leaf_61_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5373_ (.D(_0535_),
    .RN(net34),
    .CLK(clknet_leaf_51_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5374_ (.D(_0536_),
    .RN(net34),
    .CLK(clknet_leaf_52_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5375_ (.D(_0537_),
    .RN(net34),
    .CLK(clknet_leaf_52_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5376_ (.D(_0538_),
    .RN(net34),
    .CLK(clknet_leaf_52_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5377_ (.D(_0539_),
    .RN(net34),
    .CLK(clknet_leaf_25_clk),
    .Q(net18));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5378_ (.D(_0540_),
    .RN(net34),
    .CLK(clknet_leaf_26_clk),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5379_ (.D(_0541_),
    .RN(net34),
    .CLK(clknet_leaf_25_clk),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5380_ (.D(_0542_),
    .RN(net34),
    .CLK(clknet_leaf_25_clk),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5381_ (.D(_0543_),
    .RN(net34),
    .CLK(clknet_leaf_28_clk),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5382_ (.D(_0544_),
    .RN(net34),
    .CLK(clknet_leaf_28_clk),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5383_ (.D(_0545_),
    .RN(net34),
    .CLK(clknet_leaf_61_clk),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5384_ (.D(_0546_),
    .RN(net34),
    .CLK(clknet_leaf_28_clk),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5385_ (.D(_0547_),
    .RN(net34),
    .CLK(clknet_leaf_50_clk),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5386_ (.D(_0548_),
    .RN(net34),
    .CLK(clknet_leaf_50_clk),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5387_ (.D(_0549_),
    .RN(net34),
    .CLK(clknet_leaf_50_clk),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5388_ (.D(_0550_),
    .RN(net34),
    .CLK(clknet_leaf_39_clk),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5389_ (.D(_0551_),
    .RN(net34),
    .CLK(clknet_leaf_51_clk),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5390_ (.D(_0552_),
    .RN(net34),
    .CLK(clknet_leaf_48_clk),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5391_ (.D(_0553_),
    .RN(net34),
    .CLK(clknet_leaf_53_clk),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5392_ (.D(_0554_),
    .RN(net34),
    .CLK(clknet_leaf_53_clk),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5393_ (.D(_0555_),
    .RN(net34),
    .CLK(clknet_leaf_14_clk),
    .Q(net47));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5394_ (.D(_0556_),
    .RN(net34),
    .CLK(clknet_leaf_17_clk),
    .Q(net51));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5395_ (.D(_0557_),
    .RN(net34),
    .CLK(clknet_leaf_13_clk),
    .Q(net52));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _5396_ (.D(_0558_),
    .RN(net34),
    .CLK(clknet_leaf_14_clk),
    .Q(net53));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6595 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(Serial_input),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(instr[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(instr[10]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(instr[11]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(instr[12]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(instr[13]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(instr[14]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(instr[15]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(instr[1]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(instr[2]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(instr[3]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(instr[4]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(instr[5]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(instr[6]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(instr[7]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(instr[8]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(instr[9]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input18 (.I(read_data[0]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input19 (.I(read_data[10]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input20 (.I(read_data[11]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input21 (.I(read_data[12]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input22 (.I(read_data[13]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input23 (.I(read_data[14]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input24 (.I(read_data[15]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input25 (.I(read_data[1]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input26 (.I(read_data[2]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input27 (.I(read_data[3]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input28 (.I(read_data[4]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input29 (.I(read_data[5]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input30 (.I(read_data[6]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input31 (.I(read_data[7]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input32 (.I(read_data[8]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input33 (.I(read_data[9]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 input34 (.I(reset),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input35 (.I(start),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output36 (.I(net36),
    .Z(Dataw_en));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output37 (.I(net37),
    .Z(Serial_output));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output38 (.I(net38),
    .Z(data_mem_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output39 (.I(net39),
    .Z(data_mem_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output40 (.I(net40),
    .Z(data_mem_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output41 (.I(net41),
    .Z(data_mem_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output42 (.I(net42),
    .Z(data_mem_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output43 (.I(net43),
    .Z(data_mem_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output44 (.I(net44),
    .Z(data_mem_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output45 (.I(net45),
    .Z(data_mem_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output46 (.I(net46),
    .Z(hlt));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output47 (.I(net47),
    .Z(instr_mem_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output48 (.I(net48),
    .Z(instr_mem_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output49 (.I(net49),
    .Z(instr_mem_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output50 (.I(net50),
    .Z(instr_mem_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output51 (.I(net51),
    .Z(instr_mem_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output52 (.I(net52),
    .Z(instr_mem_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output53 (.I(net53),
    .Z(instr_mem_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output54 (.I(net54),
    .Z(instr_mem_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output55 (.I(net55),
    .Z(instr_mem_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output56 (.I(net56),
    .Z(instr_mem_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output57 (.I(net57),
    .Z(instr_mem_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output58 (.I(net58),
    .Z(instr_mem_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output59 (.I(net59),
    .Z(instr_mem_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output60 (.I(net60),
    .Z(write_data[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output61 (.I(net61),
    .Z(write_data[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output62 (.I(net62),
    .Z(write_data[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output63 (.I(net63),
    .Z(write_data[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output64 (.I(net64),
    .Z(write_data[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output65 (.I(net65),
    .Z(write_data[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output66 (.I(net66),
    .Z(write_data[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output67 (.I(net67),
    .Z(write_data[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output68 (.I(net68),
    .Z(write_data[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output69 (.I(net69),
    .Z(write_data[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output70 (.I(net70),
    .Z(write_data[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output71 (.I(net71),
    .Z(write_data[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output72 (.I(net72),
    .Z(write_data[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output73 (.I(net73),
    .Z(write_data[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output74 (.I(net74),
    .Z(write_data[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output75 (.I(net75),
    .Z(write_data[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_clk (.I(clknet_4_2_0_clk),
    .Z(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_clk (.I(clknet_4_2_0_clk),
    .Z(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_clk (.I(clknet_4_1_0_clk),
    .Z(clknet_leaf_2_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_clk (.I(clknet_4_3_0_clk),
    .Z(clknet_leaf_3_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_leaf_5_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_clk (.I(clknet_4_5_0_clk),
    .Z(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_clk (.I(clknet_4_5_0_clk),
    .Z(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_clk (.I(clknet_4_5_0_clk),
    .Z(clknet_leaf_10_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_clk (.I(clknet_4_5_0_clk),
    .Z(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_clk (.I(clknet_4_5_0_clk),
    .Z(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_clk (.I(clknet_4_5_0_clk),
    .Z(clknet_leaf_14_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_clk (.I(clknet_4_5_0_clk),
    .Z(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_clk (.I(clknet_4_7_0_clk),
    .Z(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_clk (.I(clknet_4_7_0_clk),
    .Z(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_clk (.I(clknet_4_4_0_clk),
    .Z(clknet_leaf_21_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_clk (.I(clknet_4_2_0_clk),
    .Z(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_clk (.I(clknet_4_2_0_clk),
    .Z(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_clk (.I(clknet_4_3_0_clk),
    .Z(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_clk (.I(clknet_4_3_0_clk),
    .Z(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_clk (.I(clknet_4_3_0_clk),
    .Z(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_clk (.I(clknet_4_3_0_clk),
    .Z(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_clk (.I(clknet_4_13_0_clk),
    .Z(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_clk (.I(clknet_4_6_0_clk),
    .Z(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_clk (.I(clknet_4_6_0_clk),
    .Z(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_clk (.I(clknet_4_6_0_clk),
    .Z(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_clk (.I(clknet_4_7_0_clk),
    .Z(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_clk (.I(clknet_4_7_0_clk),
    .Z(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_clk (.I(clknet_4_13_0_clk),
    .Z(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_clk (.I(clknet_4_13_0_clk),
    .Z(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_clk (.I(clknet_4_13_0_clk),
    .Z(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_clk (.I(clknet_4_13_0_clk),
    .Z(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_43_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_44_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_48_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_49_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_clk (.I(clknet_4_15_0_clk),
    .Z(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_56_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_leaf_62_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_leaf_63_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_clk (.I(clknet_4_2_0_clk),
    .Z(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_clk (.I(clknet_4_12_0_clk),
    .Z(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_clk (.I(clknet_4_14_0_clk),
    .Z(clknet_leaf_77_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_leaf_81_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_clk (.I(clknet_4_11_0_clk),
    .Z(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_84_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_leaf_86_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_leaf_87_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_leaf_88_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_leaf_90_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_clk (.I(clknet_4_10_0_clk),
    .Z(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_clk (.I(clknet_4_8_0_clk),
    .Z(clknet_leaf_101_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_leaf_103_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_leaf_104_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_leaf_105_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_clk (.I(clknet_4_9_0_clk),
    .Z(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_108_clk (.I(clknet_4_2_0_clk),
    .Z(clknet_leaf_108_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_109_clk (.I(clknet_4_1_0_clk),
    .Z(clknet_leaf_109_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_110_clk (.I(clknet_4_0_0_clk),
    .Z(clknet_leaf_110_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_112_clk (.I(clknet_4_0_0_clk),
    .Z(clknet_leaf_112_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_113_clk (.I(clknet_4_0_0_clk),
    .Z(clknet_leaf_113_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_114_clk (.I(clknet_4_0_0_clk),
    .Z(clknet_leaf_114_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_115_clk (.I(clknet_4_0_0_clk),
    .Z(clknet_leaf_115_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_116_clk (.I(clknet_4_0_0_clk),
    .Z(clknet_leaf_116_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_117_clk (.I(clknet_4_0_0_clk),
    .Z(clknet_leaf_117_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_118_clk (.I(clknet_4_1_0_clk),
    .Z(clknet_leaf_118_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_119_clk (.I(clknet_4_1_0_clk),
    .Z(clknet_leaf_119_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_120_clk (.I(clknet_4_1_0_clk),
    .Z(clknet_leaf_120_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_121_clk (.I(clknet_4_2_0_clk),
    .Z(clknet_leaf_121_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_clk (.I(clk),
    .Z(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_0_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_1_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_2_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_3_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_4_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_5_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_6_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_7_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_8_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_9_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_10_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_11_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_12_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_13_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_14_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_15_0_clk (.I(clknet_0_clk),
    .Z(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2639__A2 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__I (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i0 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A1 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__A2 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__I (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__B2 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A1 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__I (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__B1 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[10].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__A1 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[11].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__A2 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[11].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A1 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[11].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2652__I (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[11].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__A2 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[14].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2728__I (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[14].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A1 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[1].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__I (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[1].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__I (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[1].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__A2 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[4].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__I (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[4].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A1 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__A2 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__A1 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__I (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[5].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A1 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[6].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__A2 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[6].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__I (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[6].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__A2 (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[7].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2583__I (.I(\Arithmetic_Logic_Unit.ALU_001.Y_CY[7].i3 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__B (.I(\Arithmetic_Logic_Unit.ALU_001.p_Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2862__I (.I(\Arithmetic_Logic_Unit.ALU_001.p_Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__A2 (.I(\Arithmetic_Logic_Unit.ALU_001.p_Z ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__D (.I(\Control_unit1.instr_decoder1.A[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2823__A1 (.I(\Control_unit1.instr_decoder1.A[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__A1 (.I(\Control_unit1.instr_decoder1.A[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__I (.I(\Control_unit1.instr_decoder1.A[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__D (.I(\Control_unit1.instr_stage1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2945__A1 (.I(\Control_unit1.instr_stage1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2829__B (.I(\Control_unit1.instr_stage1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2769__A1 (.I(\Control_unit1.instr_stage1[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__D (.I(\Control_unit1.instr_stage1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2817__A1 (.I(\Control_unit1.instr_stage1[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__D (.I(\Control_unit1.instr_stage1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2826__A2 (.I(\Control_unit1.instr_stage1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2770__A2 (.I(\Control_unit1.instr_stage1[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__D (.I(\Control_unit1.instr_stage1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2826__A1 (.I(\Control_unit1.instr_stage1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2770__A1 (.I(\Control_unit1.instr_stage1[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__D (.I(\Control_unit1.instr_stage1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__A1 (.I(\Control_unit1.instr_stage1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__A1 (.I(\Control_unit1.instr_stage1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__A2 (.I(\Control_unit1.instr_stage1[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__D (.I(\Control_unit1.instr_stage1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__B2 (.I(\Control_unit1.instr_stage1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__A2 (.I(\Control_unit1.instr_stage1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__A2 (.I(\Control_unit1.instr_stage1[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__D (.I(\Control_unit1.instr_stage1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__A1 (.I(\Control_unit1.instr_stage1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__A1 (.I(\Control_unit1.instr_stage1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__A1 (.I(\Control_unit1.instr_stage1[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__D (.I(\Control_unit1.instr_stage1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__A1 (.I(\Control_unit1.instr_stage1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2789__A1 (.I(\Control_unit1.instr_stage1[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__D (.I(\Control_unit1.instr_stage1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__A1 (.I(\Control_unit1.instr_stage1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2794__A1 (.I(\Control_unit1.instr_stage1[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__D (.I(\Control_unit1.instr_stage1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__A1 (.I(\Control_unit1.instr_stage1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2800__A1 (.I(\Control_unit1.instr_stage1[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__D (.I(\Control_unit1.instr_stage1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2859__A1 (.I(\Control_unit1.instr_stage1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__A1 (.I(\Control_unit1.instr_stage1[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__D (.I(\Control_unit1.instr_stage1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__A1 (.I(\Control_unit1.instr_stage1[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__D (.I(\Control_unit1.instr_stage1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2813__A1 (.I(\Control_unit1.instr_stage1[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3083__A2 (.I(\Control_unit2.instr_decoder2.A[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__C (.I(\Control_unit2.instr_decoder2.A[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__I (.I(\Control_unit2.instr_decoder2.A[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A2 (.I(\Control_unit2.instr_decoder2.A[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__B (.I(\Control_unit2.instr_decoder2.A[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__A1 (.I(\Control_unit2.instr_decoder2.A[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__I (.I(\Control_unit2.instr_decoder2.A[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3199__I (.I(\Control_unit2.instr_stage2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__A3 (.I(\Control_unit2.instr_stage2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__A2 (.I(\Control_unit2.instr_stage2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__I (.I(\Control_unit2.instr_stage2[10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2932__I (.I(\Control_unit2.instr_stage2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__I (.I(\Control_unit2.instr_stage2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__A2 (.I(\Control_unit2.instr_stage2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__A2 (.I(\Control_unit2.instr_stage2[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A1 (.I(\Control_unit2.instr_stage2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2846__A1 (.I(\Control_unit2.instr_stage2[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2878__A1 (.I(\Control_unit2.instr_stage2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__A1 (.I(\Control_unit2.instr_stage2[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__A1 (.I(\Control_unit2.instr_stage2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2852__A1 (.I(\Control_unit2.instr_stage2[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2898__A1 (.I(\Control_unit2.instr_stage2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__A1 (.I(\Control_unit2.instr_stage2[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__A1 (.I(\Control_unit2.instr_stage2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2858__A1 (.I(\Control_unit2.instr_stage2[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__A1 (.I(\Control_unit2.instr_stage2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3150__I (.I(\Control_unit2.instr_stage2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2911__I (.I(\Control_unit2.instr_stage2[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3284__I (.I(\Control_unit2.instr_stage2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3151__A2 (.I(\Control_unit2.instr_stage2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3081__A1 (.I(\Control_unit2.instr_stage2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2917__I (.I(\Control_unit2.instr_stage2[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(Serial_input));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2825__I (.I(\Stack_pointer.SP[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2779__A1 (.I(\Stack_pointer.SP[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__A1 (.I(\Stack_pointer.SP[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2773__A1 (.I(\Stack_pointer.SP[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2840__B2 (.I(\Stack_pointer.SP[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2788__A1 (.I(\Stack_pointer.SP[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2786__A1 (.I(\Stack_pointer.SP[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2781__A1 (.I(\Stack_pointer.SP[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__C2 (.I(\Stack_pointer.SP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2793__A1 (.I(\Stack_pointer.SP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2792__A1 (.I(\Stack_pointer.SP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__A1 (.I(\Stack_pointer.SP[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__B2 (.I(\Stack_pointer.SP[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__A1 (.I(\Stack_pointer.SP[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2797__A1 (.I(\Stack_pointer.SP[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__A1 (.I(\Stack_pointer.SP[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__B2 (.I(\Stack_pointer.SP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__A1 (.I(\Stack_pointer.SP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__A1 (.I(\Stack_pointer.SP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2802__A1 (.I(\Stack_pointer.SP[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2856__B2 (.I(\Stack_pointer.SP[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2812__A1 (.I(\Stack_pointer.SP[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2811__A1 (.I(\Stack_pointer.SP[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2859__B2 (.I(\Stack_pointer.SP[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2816__A1 (.I(\Stack_pointer.SP[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2815__A1 (.I(\Stack_pointer.SP[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__D (.I(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__D (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__D (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__D (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2749__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2704__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__I1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__C2 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__A2 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__B1 (.I(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__A1 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__I (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3261__I (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__I0 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__I (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3074__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2750__A1 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__A3 (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__C (.I(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__I1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__C2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__A2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__B1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3145__A2 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__A2 (.I(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__I (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__I (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3268__I (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__I (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2755__I (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2753__A1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2752__A2 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__B1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3273__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__I (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3194__A1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3127__A1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3021__A1 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__I (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__B2 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3064__I1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__A2 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3278__I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2758__I (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2837__I (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2819__I (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A2 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__I (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__I (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__I (.I(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2815__A2 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2787__I (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2766__I (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__I (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2782__I (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__I (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2772__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2784__I (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2775__I (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2772__A2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__A1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__B2 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2922__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2836__I (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2824__I (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2828__A1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2852__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2846__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2835__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2894__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__I (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2838__A2 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__A2 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3134__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3083__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__I (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__A1 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3078__A1 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3077__B (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2844__A1 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__I (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3149__A1 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3147__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2863__B (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__C (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2883__I (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2871__I (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2944__B1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__B1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__B1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__B1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__B1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2935__B1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__I (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2944__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__A2 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__B1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__B1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2915__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2943__S (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2924__B (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__B1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__B1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3650__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3336__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3082__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2935__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__B1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__B1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__B1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2915__B1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3336__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3200__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2922__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__B2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__B (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3650__A3 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__A3 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3285__A3 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__A1 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__A2 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__A2 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__A2 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2935__A1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2952__I (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2948__I (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3008__I (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2988__I (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2970__I (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2949__I (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A1 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3289__I (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3031__A1 (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2951__I (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3208__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3159__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3092__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2954__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3011__I (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2991__I (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2973__I (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2953__I (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A1 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3294__I (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3033__A1 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2957__I (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__A1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3161__A1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3094__A1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2958__A1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3297__I (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3035__A1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2961__I (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3163__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3096__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2962__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3300__I (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3038__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2965__I (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3165__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3098__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2966__A1 (.I(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A1 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3524__I (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3303__I (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2969__I (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3226__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3170__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3103__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2975__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3223__I (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2972__I (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3169__A1 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3102__A1 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__I0 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2974__A1 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__A1 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__A1 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3229__I (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2977__I (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3171__A1 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3104__A1 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__I0 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2978__A1 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__A1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A1 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3234__I (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2981__I (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3173__A1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3106__A1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__I0 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2982__A1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__A1 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3239__I (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2985__I (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3175__A1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3108__A1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__I0 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2986__A1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A1 (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3245__I (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2990__I (.I(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3179__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3112__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__I0 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2992__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3251__I (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2995__I (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3181__A1 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3114__A1 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3051__I0 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2996__A1 (.I(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A1 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3320__I (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3053__A1 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2999__I (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3256__A1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3183__A1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3116__A1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3000__A1 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__I (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3323__I (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3003__I (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3260__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3186__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3119__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3007__A1 (.I(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3258__I (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3005__I (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3185__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3118__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3056__I0 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3006__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3264__I (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3010__I (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3122__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3058__I0 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3012__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__A1 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A1 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3270__I (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3015__I (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3124__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__I0 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3016__A1 (.I(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3275__I (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3019__I (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3126__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__I0 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3020__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3280__I (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3023__I (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__A1 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__A1 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3064__I0 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3024__A1 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3037__I (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3030__I (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3028__I (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3064__S (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3055__I (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3044__I (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3029__I (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3039__A2 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3036__A2 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3034__A2 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3032__A2 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3054__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3035__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3033__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3031__A2 (.I(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3062__S (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3060__S (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3058__S (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3056__S (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3148__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__B (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3079__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3069__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__A1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__A1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__A1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3560__A2 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3201__A2 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__A3 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3085__A3 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__I (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3086__I (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4236__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3087__A2 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3090__I (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3088__I (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3120__I (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3110__I (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3100__I (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3089__I (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3095__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3121__I (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3111__I (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3101__I (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3091__I (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3129__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3127__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3125__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3123__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3128__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3126__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3124__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3122__A2 (.I(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3135__A2 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3138__A4 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3139__A2 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3144__A2 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A1 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__A2 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__A1 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3154__A1 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3283__I (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3153__I (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3157__I (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3155__I (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3187__I (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3177__I (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3167__I (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3156__I (.I(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3188__I (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3178__I (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3168__I (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3158__I (.I(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3186__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3184__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3182__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3180__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3196__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3194__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3192__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3190__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3195__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3193__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3191__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3189__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A1 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__A1 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3423__I (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3198__I (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3386__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3343__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3293__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3209__A1 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4236__A2 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__A1 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3380__A2 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__A1 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__I (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3202__I (.I(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A2 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__A2 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3203__A2 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3206__I (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3204__I (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3263__I (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3244__I (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3222__I (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3205__I (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3265__I (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3246__I (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3224__I (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3207__I (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3220__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3216__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3212__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3208__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__A1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__I (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3211__I (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3388__A1 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3345__A1 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3296__A1 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3213__A1 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3434__I (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3215__I (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3390__A1 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3347__A1 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3299__A1 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3217__A1 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__A1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3437__I (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3219__I (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3392__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3349__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3302__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3221__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__A1 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A1 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3446__I (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3228__I (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3398__A1 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3355__A1 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3309__A1 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3231__A1 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__I (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3233__I (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__A1 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3357__A1 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3311__A1 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3236__A1 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__A1 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A1 (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3456__I (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3238__I (.I(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3402__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3359__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3313__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3241__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__A1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__I (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3243__I (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3406__A1 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3363__A1 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3317__A1 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3248__A1 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A1 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__I (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3250__I (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__A1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3365__A1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3319__A1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3253__A1 (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3410__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3367__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3322__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3257__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3368__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3324__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3259__A1 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__A1 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A1 (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3480__I (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3262__I (.I(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3282__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3277__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3272__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3267__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3281__A2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3276__A2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3271__A2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3266__A2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3487__I (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3269__I (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__A1 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A1 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3492__I (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3274__I (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3377__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3277__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__A1 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__A1 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3497__I (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3279__I (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3422__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3379__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3282__A1 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A2 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__A2 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__A1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3286__A2 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3290__I (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3287__I (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3326__I (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3314__I (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3304__I (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3288__I (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3385__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3342__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3292__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3327__I (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3315__I (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3305__I (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3291__I (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3387__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3344__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3295__A1 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3389__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3346__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3298__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3391__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3348__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3301__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3396__A1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3353__A1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3307__A1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3474__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3409__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3366__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3321__A1 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__A1 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3412__A1 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3369__A1 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3325__A1 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3335__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3333__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3331__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3329__A2 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3334__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3332__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3330__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3328__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A2 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__A2 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3337__A2 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3340__I (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3338__I (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3370__I (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3360__I (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3350__I (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3339__I (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3371__I (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3361__I (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3351__I (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3341__I (.I(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3379__A2 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3377__A2 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3375__A2 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3373__A2 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3383__I (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3381__I (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3413__I (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3403__I (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3393__I (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3382__I (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3414__I (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3404__I (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3394__I (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3384__I (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3422__A2 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__A2 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3418__A2 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3416__A2 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3417__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3415__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3568__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3481__I (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3462__I (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__I (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3426__I (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__I (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__I (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3443__I (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__I (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3515__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3615__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3572__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3519__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3436__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3574__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__I (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__I (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__I (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3442__I (.I(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3620__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3577__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3527__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__A1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__A1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3530__A1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3450__A1 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__I (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__I (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__I (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__I (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3529__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__A1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3582__A1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__A1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3455__A1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__I (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__I (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3682__I (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__I (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3584__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3534__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__I (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__I (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__I (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__I (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__A1 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3583__A1 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3533__A1 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__A1 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A1 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__A1 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3538__A1 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__A1 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__I (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__I (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__I (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__I (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3587__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3537__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3466__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__A1 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__I (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__I (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__I (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__I (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__A1 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__A1 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__A1 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__A1 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3544__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__I (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3917__I (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__I (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3477__I (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3593__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3478__A1 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3501__A2 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3496__A2 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__A2 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3486__A2 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__I (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__I (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__I (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3483__I (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__A2 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3495__A2 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3490__A2 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__A2 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__A1 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__A1 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3553__A1 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__A1 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__I (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3927__I (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3718__I (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__I (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__A1 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A1 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__A1 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3490__A1 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__I (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3931__I (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__I (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__I (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3495__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__I (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__I (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__I (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__I (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__A1 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A1 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3556__A1 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3500__A1 (.I(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__A2 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A2 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A1 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3503__A2 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3508__I (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3504__I (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__I (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3535__I (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__I (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3505__I (.I(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__I (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__I (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__I (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__I (.I(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3610__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3510__A1 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__I (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__I (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__I (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3509__I (.I(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__I (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__I (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__I (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3513__I (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3569__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3514__A1 (.I(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__I (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__I (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__I (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3517__I (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3518__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__A1 (.I(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3547__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3557__A2 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3555__A2 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3553__A2 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3551__A2 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A2 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A2 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__A2 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3562__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__I (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__I (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__A2 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__A1 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3605__A2 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3562__A2 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__I (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3585__I (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__I (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__I (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__I (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3586__I (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3576__I (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3566__I (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3638__I (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__I (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__I (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__I (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__I (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__I (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__I (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__I (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__I (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__I (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__I (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3649__I (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__A1 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__A1 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__A1 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__A1 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__I (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__I (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__I (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__I (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4288__I (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__I (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__I (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__I (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__A1 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__A1 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__A1 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3661__A1 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__I (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__I (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__I (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__I (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3793__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__I (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__I (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__I (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__I (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A1 (.I(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3842__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3798__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3752__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__A1 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__I (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4097__I (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__I (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__I (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__I (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__I (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__I (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__I (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__I (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__I (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__I (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3686__I (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4314__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3691__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__A2 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__A2 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A2 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__A2 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__I (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__I (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__I (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3698__I (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__I (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__I (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__I (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__I (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__I (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__I (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__I (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__I (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3725__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3715__A2 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__I (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__I (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__I (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__I (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__A1 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__A1 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__A1 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__A1 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4340__I (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__I (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__I (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__I (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__I (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4139__I (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__I (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__I (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__I (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__I (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__I (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__I (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3788__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__I (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__I (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__I (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3736__I (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__A1 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A1 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__A1 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3740__A1 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__I (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__I (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__I (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__I (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3799__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3753__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__A2 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__A2 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__A2 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3763__A2 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__A1 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__A1 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__A1 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__A1 (.I(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__I (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__I (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__I (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__I (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3919__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__A2 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__A2 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__A2 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__A2 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__I (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__I (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__I (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__I (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__I (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__I (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__I (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3787__I (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__A2 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__A2 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__A2 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__A2 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__A2 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__A2 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3820__A2 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__A2 (.I(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A2 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A2 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A2 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__A2 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__I (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__I (.I(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__I (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__I (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__I (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__I (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__A2 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A2 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A2 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__A2 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A2 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__A2 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__A2 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__A2 (.I(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A1 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__A1 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A1 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A1 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__I (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__I (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__I (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__I (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__I (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__I (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A2 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A2 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A2 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A2 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__I (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3907__I (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__I (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__I (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__A1 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A1 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__A1 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A1 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A2 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__A2 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__A2 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__A2 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3902__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__A2 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__A2 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3912__A2 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__A2 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3925__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__A2 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3932__A2 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__A2 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__A2 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__I (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__I (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__I (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__I (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__I (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__I (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A2 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A2 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__A2 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A2 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__A1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__A1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__A1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__I (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3967__I (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__I (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__I (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__A1 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A1 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__A1 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__A1 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__A2 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__A2 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__A2 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__A2 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3964__A2 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__A2 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3960__A2 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__A2 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__A2 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A2 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A2 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3981__A2 (.I(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A2 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__A2 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A2 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A2 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__I (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__I (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__I (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__I (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__I (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__I (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A2 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__A2 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A2 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__A2 (.I(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A2 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__A2 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__A2 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__A2 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__A2 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__A2 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__A2 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__A2 (.I(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__A2 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__A2 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__A2 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A2 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__A2 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__A2 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__A2 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__A2 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__A2 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A2 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__A2 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A2 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__I (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__I (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__I (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__I (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__I (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__I (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A2 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A2 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__A2 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A2 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__I (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__I (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__I (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__I (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A2 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A2 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A2 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A2 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__A2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__A2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A2 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__A2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4051__A2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__A2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A2 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A2 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A2 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__A2 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__A2 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__A2 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__A2 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__A2 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4073__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__I (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__I (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__I (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__I (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__I (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__I (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__I (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4112__I (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__I (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__I (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4090__A2 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A2 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A2 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__A2 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4244__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__A1 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__A1 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__A1 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__A1 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A1 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4181__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A2 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A2 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A2 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4130__A2 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__A1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__A1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__A1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__A2 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__A2 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A2 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__A2 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__A1 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__A1 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__A1 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A1 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4275__A1 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4232__A1 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__A1 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4137__A1 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__I (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__I (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__I (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__I (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4161__I (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__I (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__A2 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__A2 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A2 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A2 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__I (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__I (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4162__I (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__I (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__A2 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4168__A2 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A2 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A2 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A2 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A2 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__A2 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__A2 (.I(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__A1 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__A1 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A1 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4178__A1 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__A1 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__A1 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__A1 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__A1 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4188__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__A2 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__A2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__A2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__A2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__A2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__I (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__I (.I(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4226__I (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4216__I (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4206__I (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4195__I (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4203__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A2 (.I(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__I (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4217__I (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__I (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__I (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4215__A2 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__A2 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4211__A2 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__A2 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__A2 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4223__A2 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__A2 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__A2 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__A2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__A2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4229__A2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4232__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__A2 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4239__I (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__I (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__I (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__I (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__I (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__I (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4248__A2 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__A2 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4244__A2 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A2 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__I (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4260__I (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__I (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__I (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__A2 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__A2 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__A2 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A2 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4256__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__A2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__A2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__A2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__A2 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__A2 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__A2 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4262__A2 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4272__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4275__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__A1 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A1 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A1 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__A1 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A1 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__A1 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A1 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A1 (.I(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4331__I (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__I (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__I (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__I (.I(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A2 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A2 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__A2 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__A2 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__I (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__I (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4299__I (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__I (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A1 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A1 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A1 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__A1 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__A1 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__A1 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__A1 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A1 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4328__A1 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4343__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__A2 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__I (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__I (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__I (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__I (.I(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__A2 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4361__A2 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A2 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A2 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__I (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__I (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__I (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__I (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__A2 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__A2 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__A2 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__A2 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__A1 (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A1 (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__A1 (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__A1 (.I(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A1 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__A1 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A1 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__A1 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A2 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__A2 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__A2 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__A2 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A2 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__A2 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A2 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A2 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__A1 (.I(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A2 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A2 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A2 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__A2 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__A2 (.I(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4411__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__I (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__I (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__I (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__I (.I(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A2 (.I(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A2 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__A2 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A2 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__A2 (.I(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A2 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__A2 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__A2 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__A2 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__A2 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__A2 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A2 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__A2 (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__A2 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__I (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__I (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__I (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__I (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4453__A2 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4451__A2 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A2 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__A2 (.I(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__I (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__I (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__I (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__I (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__A2 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__A2 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A2 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A2 (.I(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__A2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4471__A2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A2 (.I(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__A2 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A2 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__A2 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A2 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A1 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A1 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A1 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A1 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4535__I (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__I (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__I (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__I (.I(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__I (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__I (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__I (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__I (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A2 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A2 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__A2 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__A2 (.I(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A1 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A1 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__A1 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__A1 (.I(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__A1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A1 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__A1 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A1 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__A1 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4500__A1 (.I(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A1 (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A1 (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__A1 (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__A1 (.I(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__A1 (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__A1 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A1 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__A1 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__A1 (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__A1 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A1 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A1 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__A1 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A1 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A1 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A1 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4523__A1 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A1 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A1 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__A1 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__A1 (.I(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A1 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__A1 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__A1 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__A1 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A2 (.I(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4550__A2 (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A2 (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A2 (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A2 (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__I (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__I (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__I (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4554__I (.I(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__A2 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A2 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__A2 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A2 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__A1 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A1 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__A1 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A1 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__I (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__I (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__I (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__I (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__A1 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A1 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A1 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A1 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A1 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__A1 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__A1 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A1 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A1 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A1 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A1 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A1 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A1 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__A1 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A1 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__A1 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A2 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__A2 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__A2 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A2 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A2 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A2 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__A2 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A2 (.I(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__I (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__I (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__I (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__I (.I(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A2 (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__A2 (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A2 (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A2 (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__I (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__I (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__I (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__I (.I(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A2 (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__A2 (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A2 (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__A2 (.I(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A2 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__A2 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A2 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__A2 (.I(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__I (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__I (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__I (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__I (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__I (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__I (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__I (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__I (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A2 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__A2 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A2 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A2 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__A2 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A2 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A2 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A2 (.I(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__A2 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A2 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__A2 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A2 (.I(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__I (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__I (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__I (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__I (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__I (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__I (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__I (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__I (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__I (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__I (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__I (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__I (.I(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__I (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__I (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__I (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__I (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__A2 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__A2 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A2 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__A2 (.I(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__A1 (.I(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A1 (.I(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__A1 (.I(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A1 (.I(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__I (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A2 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2832__A1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2432__A1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2424__I (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__A1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__A1 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__A1 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__A1 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2387__I (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__A1 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__A1 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__A1 (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2388__I (.I(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A1 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__A1 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2835__A1 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A3 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2830__A2 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__A1 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A4 (.I(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3152__A1 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2942__A1 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__A1 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__A1 (.I(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2412__I (.I(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__I (.I(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2574__A2 (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__A2 (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__I (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__I (.I(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__B2 (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__B2 (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__B (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2405__B (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2525__A3 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A3 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A4 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2410__A4 (.I(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3068__A1 (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__C2 (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__A2 (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__A1 (.I(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A2 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__I (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2525__A2 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2417__A2 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A2 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__I (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2415__I (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__S (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__S (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__B2 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__C2 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__A2 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__B2 (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3084__A1 (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__B (.I(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__A1 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__A1 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__A1 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__A1 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2639__A1 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__A1 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__A2 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2534__A2 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2524__A2 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__A2 (.I(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2575__A1 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__A1 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__A1 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__I (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2716__A1 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__A1 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__A1 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2437__I (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__A2 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__C2 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__A2 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__B1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__A2 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A2 (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2472__I (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__I (.I(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__B1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__B1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__I (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__I (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3146__A1 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__I1 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3083__B (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__A1 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2453__I (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__I (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__A1 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2540__A1 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2468__I (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__I (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__S (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2569__I (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__I (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__S (.I(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__A1 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__I (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3197__I (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__I (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3160__A1 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3093__A1 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2955__A1 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2452__I (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2686__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2591__I (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__I (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2709__A1 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__A1 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__A1 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A1 (.I(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__B1 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A3 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A3 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__A3 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__I (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__B2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__B2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__B (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__A1 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__C (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__A2 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2464__A1 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__I (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2576__A2 (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2530__A2 (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2462__A2 (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__A2 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2482__A3 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2464__A2 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__A3 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__C2 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A2 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2474__B1 (.I(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__A2 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A1 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__I (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3210__I (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__I (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3162__A1 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3095__A1 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2959__A1 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__I (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__A2 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__A2 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A1 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__A1 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A1 (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__I (.I(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3141__A4 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__B2 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A2 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__B1 (.I(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__A2 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A1 (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__I (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3214__I (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__I (.I(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3164__A1 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3097__A1 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2963__A1 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__I (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A2 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__A2 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A2 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__A2 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2526__A2 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__A3 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2506__A1 (.I(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__A2 (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2527__A2 (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__A4 (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2506__A2 (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3137__A1 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__I0 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__A1 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3040__I1 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__B2 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__B1 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2756__B1 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__B2 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__B2 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__B2 (.I(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__C1 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__C1 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__C1 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__C1 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__I1 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A1 (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__I (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3218__I (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__I (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3166__A1 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3099__A1 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2967__A1 (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__I (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__A1 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__I (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2573__A1 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A1 (.I(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__B (.I(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__I (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__I (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2968__I (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2542__I (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3147__C (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3067__I (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3066__A2 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__A1 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2657__I (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__A2 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2603__A2 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__A2 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__S (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2745__S (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__A1 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__A1 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__A3 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3045__I1 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2898__B2 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A1 (.I(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__B1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__C1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__C1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__I (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__B (.I(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__I (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__I (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3227__I (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__I (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__A2 (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__A2 (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2698__A2 (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__I (.I(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3075__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2751__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2715__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2573__A2 (.I(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__A1 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A1 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2598__A1 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__I (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3047__I1 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__B2 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__C2 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__A1 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3140__A2 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3042__I1 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__B2 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__B2 (.I(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__A3 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__B (.I(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__I (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__I (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3232__I (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__I (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__B (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__B (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__A1 (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__B1 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__A1 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__C2 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A1 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__A1 (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2595__I (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3049__I1 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__B2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__A1 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3144__A1 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__A2 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3137__A2 (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2608__A2 (.I(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__I (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__I (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3237__I (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__I (.I(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3132__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2623__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A3 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A2 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2622__A2 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3131__A1 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2702__A1 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A1 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2628__A1 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3051__I1 (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__B2 (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__A2 (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__B1 (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3143__A1 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__A2 (.I(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4518__I (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__I (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3242__I (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2635__I (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3143__A2 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__I1 (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__I (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3249__I (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__A1 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2650__I (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3182__A1 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3115__A1 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2997__A1 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2651__I (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3056__I1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__C2 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2698__A1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__A1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A3 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__C (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2924__A1 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A1 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__A2 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2718__A2 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__A2 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__A2 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__A2 (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__A2 (.I(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2924__A2 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A2 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__I (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__I (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3254__I (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2670__I (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3058__I1 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__C2 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2708__A2 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__A1 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2686__B (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__I (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3769__I (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3002__I (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__I (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2714__A1 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__A2 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_clk_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(instr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(instr[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(instr[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(instr[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(instr[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(instr[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(instr[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(instr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(instr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(instr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(instr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(instr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(instr[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(instr[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(instr[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(instr[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(read_data[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(read_data[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(read_data[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(read_data[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(read_data[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(read_data[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(read_data[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(read_data[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(read_data[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(read_data[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(read_data[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(read_data[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(read_data[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(read_data[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(read_data[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(read_data[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(reset));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(start));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2427__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__I1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__D (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__D (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__D (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__D (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__D (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__D (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2950__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2998__I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3476__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3004__I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3482__I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3009__I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3488__I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3014__I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3018__I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3022__I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4356__I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3512__I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2956__I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4359__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3516__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2960__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4362__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3520__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2964__I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4298__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2971__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4507__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2976__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4307__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2980__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2984__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3463__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2989__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4321__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2994__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__SETN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__SETN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__SETN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__SETN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__RN (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2879__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__B (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__I0 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output41_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output42_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output43_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output44_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output45_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output46_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2879__A2 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output47_I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__A1 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output48_I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2926__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output49_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2939__A1 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2936__I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2934__A1 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output50_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2940__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output51_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__A2 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A2 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__A2 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output52_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A3 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__A3 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output53_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__A4 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output54_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2884__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output55_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__A1 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2890__I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2886__A1 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__A1 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output56_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__A2 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2896__A1 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2892__I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output57_I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2902__A1 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output58_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2907__A1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output59_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__A2 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__A1 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output60_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output61_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output62_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__A1 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output63_I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output64_I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output65_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output66_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output67_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output68_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output69_I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output70_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output71_I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output72_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output73_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output74_I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output75_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__CLK (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__CLK (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__CLK (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__CLK (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__CLK (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__CLK (.I(clknet_leaf_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__CLK (.I(clknet_leaf_1_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__CLK (.I(clknet_leaf_4_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__CLK (.I(clknet_leaf_6_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__CLK (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4798__CLK (.I(clknet_leaf_7_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__CLK (.I(clknet_leaf_8_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__CLK (.I(clknet_leaf_11_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__CLK (.I(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__CLK (.I(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__CLK (.I(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__CLK (.I(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__CLK (.I(clknet_leaf_12_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__CLK (.I(clknet_leaf_13_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__CLK (.I(clknet_leaf_15_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__CLK (.I(clknet_leaf_17_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__CLK (.I(clknet_leaf_18_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__CLK (.I(clknet_leaf_19_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__CLK (.I(clknet_leaf_22_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__CLK (.I(clknet_leaf_23_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__CLK (.I(clknet_leaf_24_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__CLK (.I(clknet_leaf_25_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__CLK (.I(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__CLK (.I(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__CLK (.I(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__CLK (.I(clknet_leaf_26_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__CLK (.I(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__CLK (.I(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__CLK (.I(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__CLK (.I(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__CLK (.I(clknet_leaf_27_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__CLK (.I(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__CLK (.I(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__CLK (.I(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__CLK (.I(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__CLK (.I(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__CLK (.I(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__CLK (.I(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__CLK (.I(clknet_leaf_28_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__CLK (.I(clknet_leaf_30_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__CLK (.I(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__CLK (.I(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4834__CLK (.I(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__CLK (.I(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__CLK (.I(clknet_leaf_31_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__CLK (.I(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__CLK (.I(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__CLK (.I(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__CLK (.I(clknet_leaf_32_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4841__CLK (.I(clknet_leaf_33_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__CLK (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__CLK (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__CLK (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__CLK (.I(clknet_leaf_34_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__CLK (.I(clknet_leaf_36_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__CLK (.I(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__CLK (.I(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__CLK (.I(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__CLK (.I(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__CLK (.I(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__CLK (.I(clknet_leaf_37_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__CLK (.I(clknet_leaf_38_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__CLK (.I(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__CLK (.I(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__CLK (.I(clknet_leaf_39_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__CLK (.I(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__CLK (.I(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4923__CLK (.I(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__CLK (.I(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__CLK (.I(clknet_leaf_40_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__CLK (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__CLK (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__CLK (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__CLK (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__CLK (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__CLK (.I(clknet_leaf_41_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__CLK (.I(clknet_leaf_42_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__CLK (.I(clknet_leaf_44_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__CLK (.I(clknet_leaf_44_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__CLK (.I(clknet_leaf_44_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__CLK (.I(clknet_leaf_44_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__CLK (.I(clknet_leaf_44_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__CLK (.I(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__CLK (.I(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__CLK (.I(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__CLK (.I(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__CLK (.I(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__CLK (.I(clknet_leaf_45_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__CLK (.I(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__CLK (.I(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__CLK (.I(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__CLK (.I(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__CLK (.I(clknet_leaf_46_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__CLK (.I(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__CLK (.I(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__CLK (.I(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__CLK (.I(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__CLK (.I(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__CLK (.I(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__CLK (.I(clknet_leaf_47_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__CLK (.I(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__CLK (.I(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__CLK (.I(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__CLK (.I(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__CLK (.I(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__CLK (.I(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__CLK (.I(clknet_leaf_50_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__CLK (.I(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__CLK (.I(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__CLK (.I(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__CLK (.I(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__CLK (.I(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__CLK (.I(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__CLK (.I(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__CLK (.I(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__CLK (.I(clknet_leaf_51_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__CLK (.I(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__CLK (.I(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__CLK (.I(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__CLK (.I(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__CLK (.I(clknet_leaf_52_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__CLK (.I(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__CLK (.I(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__CLK (.I(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__CLK (.I(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__CLK (.I(clknet_leaf_53_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5312__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__CLK (.I(clknet_leaf_54_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__CLK (.I(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__CLK (.I(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__CLK (.I(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__CLK (.I(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__CLK (.I(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__CLK (.I(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__CLK (.I(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__CLK (.I(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__CLK (.I(clknet_leaf_55_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__CLK (.I(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__CLK (.I(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__CLK (.I(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__CLK (.I(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__CLK (.I(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__CLK (.I(clknet_leaf_57_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__CLK (.I(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__CLK (.I(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__CLK (.I(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__CLK (.I(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__CLK (.I(clknet_leaf_58_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__CLK (.I(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__CLK (.I(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__CLK (.I(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__CLK (.I(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__CLK (.I(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__CLK (.I(clknet_leaf_59_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__CLK (.I(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__CLK (.I(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__CLK (.I(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__CLK (.I(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__CLK (.I(clknet_leaf_60_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__CLK (.I(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__CLK (.I(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__CLK (.I(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__CLK (.I(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__CLK (.I(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__CLK (.I(clknet_leaf_61_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__CLK (.I(clknet_leaf_62_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__CLK (.I(clknet_leaf_62_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__CLK (.I(clknet_leaf_62_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__CLK (.I(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__CLK (.I(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__CLK (.I(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__CLK (.I(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__CLK (.I(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__CLK (.I(clknet_leaf_64_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__CLK (.I(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__CLK (.I(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__CLK (.I(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__CLK (.I(clknet_leaf_65_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__CLK (.I(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__CLK (.I(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__CLK (.I(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__CLK (.I(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__CLK (.I(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__CLK (.I(clknet_leaf_66_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__CLK (.I(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__CLK (.I(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__CLK (.I(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__CLK (.I(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5302__CLK (.I(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__CLK (.I(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__CLK (.I(clknet_leaf_67_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__CLK (.I(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__CLK (.I(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__CLK (.I(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__CLK (.I(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__CLK (.I(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__CLK (.I(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__CLK (.I(clknet_leaf_68_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__CLK (.I(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__CLK (.I(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__CLK (.I(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__CLK (.I(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__CLK (.I(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__CLK (.I(clknet_leaf_69_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__CLK (.I(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__CLK (.I(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__CLK (.I(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__CLK (.I(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__CLK (.I(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__CLK (.I(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__CLK (.I(clknet_leaf_70_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__CLK (.I(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__CLK (.I(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__CLK (.I(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__CLK (.I(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__CLK (.I(clknet_leaf_71_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__CLK (.I(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__CLK (.I(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__CLK (.I(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__CLK (.I(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__CLK (.I(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__CLK (.I(clknet_leaf_72_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__CLK (.I(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__CLK (.I(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__CLK (.I(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__CLK (.I(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__CLK (.I(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__CLK (.I(clknet_leaf_73_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__CLK (.I(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__CLK (.I(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__CLK (.I(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__CLK (.I(clknet_leaf_74_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__CLK (.I(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__CLK (.I(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__CLK (.I(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__CLK (.I(clknet_leaf_75_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__CLK (.I(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__CLK (.I(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__CLK (.I(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__CLK (.I(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__CLK (.I(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__CLK (.I(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__CLK (.I(clknet_leaf_76_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__CLK (.I(clknet_leaf_77_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__CLK (.I(clknet_leaf_77_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__CLK (.I(clknet_leaf_77_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__CLK (.I(clknet_leaf_77_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__CLK (.I(clknet_leaf_77_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__CLK (.I(clknet_leaf_77_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__CLK (.I(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__CLK (.I(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__CLK (.I(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__CLK (.I(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__CLK (.I(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__CLK (.I(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__CLK (.I(clknet_leaf_78_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__CLK (.I(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__CLK (.I(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__CLK (.I(clknet_leaf_79_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__CLK (.I(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__CLK (.I(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__CLK (.I(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__CLK (.I(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__CLK (.I(clknet_leaf_80_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__CLK (.I(clknet_leaf_81_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__CLK (.I(clknet_leaf_81_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__CLK (.I(clknet_leaf_81_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__CLK (.I(clknet_leaf_81_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__CLK (.I(clknet_leaf_81_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__CLK (.I(clknet_leaf_81_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__CLK (.I(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__CLK (.I(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__CLK (.I(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__CLK (.I(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__CLK (.I(clknet_leaf_82_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__CLK (.I(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__CLK (.I(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__CLK (.I(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__CLK (.I(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__CLK (.I(clknet_leaf_83_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__CLK (.I(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__CLK (.I(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__CLK (.I(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__CLK (.I(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__CLK (.I(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__CLK (.I(clknet_leaf_84_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__CLK (.I(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__CLK (.I(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__CLK (.I(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__CLK (.I(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__CLK (.I(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__CLK (.I(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__CLK (.I(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__CLK (.I(clknet_leaf_85_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__CLK (.I(clknet_leaf_86_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__CLK (.I(clknet_leaf_86_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__CLK (.I(clknet_leaf_86_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__CLK (.I(clknet_leaf_86_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__CLK (.I(clknet_leaf_86_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__CLK (.I(clknet_leaf_86_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__CLK (.I(clknet_leaf_87_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__CLK (.I(clknet_leaf_87_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__CLK (.I(clknet_leaf_87_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__CLK (.I(clknet_leaf_87_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__CLK (.I(clknet_leaf_87_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__CLK (.I(clknet_leaf_87_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__CLK (.I(clknet_leaf_87_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__CLK (.I(clknet_leaf_87_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__CLK (.I(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__CLK (.I(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__CLK (.I(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__CLK (.I(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__CLK (.I(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__CLK (.I(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__CLK (.I(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__CLK (.I(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__CLK (.I(clknet_leaf_91_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__CLK (.I(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__CLK (.I(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__CLK (.I(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__CLK (.I(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__CLK (.I(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__CLK (.I(clknet_leaf_92_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__CLK (.I(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__CLK (.I(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__CLK (.I(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__CLK (.I(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__CLK (.I(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__CLK (.I(clknet_leaf_93_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__CLK (.I(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__CLK (.I(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__CLK (.I(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__CLK (.I(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__CLK (.I(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__CLK (.I(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__CLK (.I(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__CLK (.I(clknet_leaf_94_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__CLK (.I(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__CLK (.I(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__CLK (.I(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__CLK (.I(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__CLK (.I(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__CLK (.I(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__CLK (.I(clknet_leaf_96_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__CLK (.I(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__CLK (.I(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__CLK (.I(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__CLK (.I(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__CLK (.I(clknet_leaf_97_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__CLK (.I(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__CLK (.I(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__CLK (.I(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__CLK (.I(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__CLK (.I(clknet_leaf_98_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__CLK (.I(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__CLK (.I(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__CLK (.I(clknet_leaf_99_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__CLK (.I(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__CLK (.I(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__CLK (.I(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__CLK (.I(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__CLK (.I(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__CLK (.I(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__CLK (.I(clknet_leaf_100_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__CLK (.I(clknet_leaf_101_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__CLK (.I(clknet_leaf_101_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__CLK (.I(clknet_leaf_101_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__CLK (.I(clknet_leaf_101_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__CLK (.I(clknet_leaf_101_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__CLK (.I(clknet_leaf_101_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__CLK (.I(clknet_leaf_101_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__CLK (.I(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__CLK (.I(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__CLK (.I(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__CLK (.I(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__CLK (.I(clknet_leaf_102_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__CLK (.I(clknet_leaf_104_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__CLK (.I(clknet_leaf_104_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__CLK (.I(clknet_leaf_104_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__CLK (.I(clknet_leaf_104_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__CLK (.I(clknet_leaf_105_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__CLK (.I(clknet_leaf_105_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__CLK (.I(clknet_leaf_105_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__CLK (.I(clknet_leaf_105_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__CLK (.I(clknet_leaf_105_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__CLK (.I(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__CLK (.I(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__CLK (.I(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__CLK (.I(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__CLK (.I(clknet_leaf_106_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__CLK (.I(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__CLK (.I(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__CLK (.I(clknet_leaf_107_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__CLK (.I(clknet_leaf_108_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__CLK (.I(clknet_leaf_108_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__CLK (.I(clknet_leaf_108_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__CLK (.I(clknet_leaf_109_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__CLK (.I(clknet_leaf_109_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__CLK (.I(clknet_leaf_109_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__CLK (.I(clknet_leaf_109_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__CLK (.I(clknet_leaf_110_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__CLK (.I(clknet_leaf_110_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__CLK (.I(clknet_leaf_110_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__CLK (.I(clknet_leaf_110_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__CLK (.I(clknet_leaf_110_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__CLK (.I(clknet_leaf_112_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__CLK (.I(clknet_leaf_112_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__CLK (.I(clknet_leaf_112_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__CLK (.I(clknet_leaf_112_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__CLK (.I(clknet_leaf_113_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__CLK (.I(clknet_leaf_113_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__CLK (.I(clknet_leaf_113_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__CLK (.I(clknet_leaf_113_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__CLK (.I(clknet_leaf_113_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__CLK (.I(clknet_leaf_113_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__CLK (.I(clknet_leaf_113_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__CLK (.I(clknet_leaf_114_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__CLK (.I(clknet_leaf_114_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__CLK (.I(clknet_leaf_114_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__CLK (.I(clknet_leaf_114_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__CLK (.I(clknet_leaf_114_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__CLK (.I(clknet_leaf_114_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__CLK (.I(clknet_leaf_114_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__CLK (.I(clknet_leaf_115_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__CLK (.I(clknet_leaf_115_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__CLK (.I(clknet_leaf_115_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__CLK (.I(clknet_leaf_115_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__CLK (.I(clknet_leaf_115_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__CLK (.I(clknet_leaf_116_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__CLK (.I(clknet_leaf_116_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__CLK (.I(clknet_leaf_116_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__CLK (.I(clknet_leaf_116_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__CLK (.I(clknet_leaf_118_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__CLK (.I(clknet_leaf_118_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__CLK (.I(clknet_leaf_118_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__CLK (.I(clknet_leaf_118_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__CLK (.I(clknet_leaf_120_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__CLK (.I(clknet_leaf_120_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__CLK (.I(clknet_leaf_120_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__CLK (.I(clknet_leaf_120_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__CLK (.I(clknet_leaf_120_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__CLK (.I(clknet_leaf_121_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__CLK (.I(clknet_leaf_121_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__CLK (.I(clknet_leaf_121_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_15_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_14_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_13_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_12_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_11_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_10_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_9_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_8_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_7_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_6_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_5_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_4_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_3_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_2_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_1_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_0_0_clk_I (.I(clknet_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_117_clk_I (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_116_clk_I (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_115_clk_I (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_114_clk_I (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_113_clk_I (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_112_clk_I (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__CLK (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_110_clk_I (.I(clknet_4_0_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_120_clk_I (.I(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_119_clk_I (.I(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_118_clk_I (.I(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_109_clk_I (.I(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_clk_I (.I(clknet_4_1_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_121_clk_I (.I(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_108_clk_I (.I(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_clk_I (.I(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_clk_I (.I(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_clk_I (.I(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_clk_I (.I(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_clk_I (.I(clknet_4_2_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_clk_I (.I(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_clk_I (.I(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_clk_I (.I(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_clk_I (.I(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_clk_I (.I(clknet_4_3_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_clk_I (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_clk_I (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_clk_I (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_clk_I (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_clk_I (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_clk_I (.I(clknet_4_4_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_clk_I (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_clk_I (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_clk_I (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_clk_I (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_clk_I (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4856__CLK (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_clk_I (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_clk_I (.I(clknet_4_5_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_clk_I (.I(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_clk_I (.I(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_clk_I (.I(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__CLK (.I(clknet_4_6_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__CLK (.I(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_clk_I (.I(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_clk_I (.I(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__CLK (.I(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_clk_I (.I(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_clk_I (.I(clknet_4_7_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_101_clk_I (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_100_clk_I (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_99_clk_I (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_98_clk_I (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_97_clk_I (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_96_clk_I (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__CLK (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_94_clk_I (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_93_clk_I (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_92_clk_I (.I(clknet_4_8_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_107_clk_I (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_106_clk_I (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_105_clk_I (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_104_clk_I (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_103_clk_I (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_102_clk_I (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_clk_I (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_clk_I (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_clk_I (.I(clknet_4_9_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_clk_I (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_90_clk_I (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__CLK (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_88_clk_I (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_87_clk_I (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_clk_I (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_clk_I (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_84_clk_I (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_83_clk_I (.I(clknet_4_10_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_clk_I (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_clk_I (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_clk_I (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_clk_I (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_clk_I (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_clk_I (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_clk_I (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_clk_I (.I(clknet_4_11_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_clk_I (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_clk_I (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_clk_I (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_clk_I (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_clk_I (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_clk_I (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_clk_I (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_clk_I (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_clk_I (.I(clknet_4_12_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_clk_I (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_clk_I (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_clk_I (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_clk_I (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__CLK (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_clk_I (.I(clknet_4_13_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_clk_I (.I(clknet_4_14_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_clk_I (.I(clknet_4_15_0_clk));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_185_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_185_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_195_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_195_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_196_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_198_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_199_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_199_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_200_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_201_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_201_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_201_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_201_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_202_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_203_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_203_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_203_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_203_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_203_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_203_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_204_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_205_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_205_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_205_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_205_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_206_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_207_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_207_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_207_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_207_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_207_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_208_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_209_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_209_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_210_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_210_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_211_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_211_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_212_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_213_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_213_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_214_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_215_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_215_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_215_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_215_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_215_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_215_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_216_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_217_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_217_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_218_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_219_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_219_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_220_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_221_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_221_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_222_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_222_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_222_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_222_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_223_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_223_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_223_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_223_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_224_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_225_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_225_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_225_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_225_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_225_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_226_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_227_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_227_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_228_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_229_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_229_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_229_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_229_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_230_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_230_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_230_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_230_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_230_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_230_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_230_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_231_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_231_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_232_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_233_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_233_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_234_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_235_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_235_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_235_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_235_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_235_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_236_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_237_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_237_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_238_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_239_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_239_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_240_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_240_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_240_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_240_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_240_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_241_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_241_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_242_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_242_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_243_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_243_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_243_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_243_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_244_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_244_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1758 ();
endmodule

