VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO io_interface
  CLASS BLOCK ;
  FOREIGN io_interface ;
  ORIGIN 0.000 0.000 ;
  SIZE 1800.000 BY 1000.000 ;
  PIN Serial_input
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1724.800 996.000 1725.360 1000.000 ;
    END
  END Serial_input
  PIN Serial_output
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1730.960 996.000 1731.520 1000.000 ;
    END
  END Serial_output
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1665.440 0.000 1666.000 4.000 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1699.040 0.000 1699.600 4.000 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1702.400 0.000 1702.960 4.000 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1705.760 0.000 1706.320 4.000 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1709.120 0.000 1709.680 4.000 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1712.480 0.000 1713.040 4.000 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1715.840 0.000 1716.400 4.000 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1719.200 0.000 1719.760 4.000 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1722.560 0.000 1723.120 4.000 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1725.920 0.000 1726.480 4.000 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1729.280 0.000 1729.840 4.000 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1668.800 0.000 1669.360 4.000 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1732.640 0.000 1733.200 4.000 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1736.000 0.000 1736.560 4.000 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1739.360 0.000 1739.920 4.000 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1742.720 0.000 1743.280 4.000 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1746.080 0.000 1746.640 4.000 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1749.440 0.000 1750.000 4.000 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1752.800 0.000 1753.360 4.000 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1756.160 0.000 1756.720 4.000 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1759.520 0.000 1760.080 4.000 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1672.160 0.000 1672.720 4.000 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1675.520 0.000 1676.080 4.000 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1678.880 0.000 1679.440 4.000 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1682.240 0.000 1682.800 4.000 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1685.600 0.000 1686.160 4.000 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1688.960 0.000 1689.520 4.000 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1692.320 0.000 1692.880 4.000 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1695.680 0.000 1696.240 4.000 ;
    END
  END analog_io[9]
  PIN clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1772.960 0.000 1773.520 4.000 ;
    END
  END clk
  PIN data_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1114.960 996.000 1115.520 1000.000 ;
    END
  END data_mem_addr[0]
  PIN data_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1139.600 996.000 1140.160 1000.000 ;
    END
  END data_mem_addr[1]
  PIN data_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1164.240 996.000 1164.800 1000.000 ;
    END
  END data_mem_addr[2]
  PIN data_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1188.880 996.000 1189.440 1000.000 ;
    END
  END data_mem_addr[3]
  PIN data_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1213.520 996.000 1214.080 1000.000 ;
    END
  END data_mem_addr[4]
  PIN data_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1238.160 996.000 1238.720 1000.000 ;
    END
  END data_mem_addr[5]
  PIN data_mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1262.800 996.000 1263.360 1000.000 ;
    END
  END data_mem_addr[6]
  PIN data_mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1287.440 996.000 1288.000 1000.000 ;
    END
  END data_mem_addr[7]
  PIN data_mem_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1102.640 996.000 1103.200 1000.000 ;
    END
  END data_mem_sel
  PIN data_read_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1121.120 996.000 1121.680 1000.000 ;
    END
  END data_read_data[0]
  PIN data_read_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1336.720 996.000 1337.280 1000.000 ;
    END
  END data_read_data[10]
  PIN data_read_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1349.040 996.000 1349.600 1000.000 ;
    END
  END data_read_data[11]
  PIN data_read_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1361.360 996.000 1361.920 1000.000 ;
    END
  END data_read_data[12]
  PIN data_read_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1373.680 996.000 1374.240 1000.000 ;
    END
  END data_read_data[13]
  PIN data_read_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1386.000 996.000 1386.560 1000.000 ;
    END
  END data_read_data[14]
  PIN data_read_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1398.320 996.000 1398.880 1000.000 ;
    END
  END data_read_data[15]
  PIN data_read_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1145.760 996.000 1146.320 1000.000 ;
    END
  END data_read_data[1]
  PIN data_read_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1170.400 996.000 1170.960 1000.000 ;
    END
  END data_read_data[2]
  PIN data_read_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1195.040 996.000 1195.600 1000.000 ;
    END
  END data_read_data[3]
  PIN data_read_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1219.680 996.000 1220.240 1000.000 ;
    END
  END data_read_data[4]
  PIN data_read_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1244.320 996.000 1244.880 1000.000 ;
    END
  END data_read_data[5]
  PIN data_read_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1268.960 996.000 1269.520 1000.000 ;
    END
  END data_read_data[6]
  PIN data_read_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1293.600 996.000 1294.160 1000.000 ;
    END
  END data_read_data[7]
  PIN data_read_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1312.080 996.000 1312.640 1000.000 ;
    END
  END data_read_data[8]
  PIN data_read_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1324.400 996.000 1324.960 1000.000 ;
    END
  END data_read_data[9]
  PIN data_write_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1127.280 996.000 1127.840 1000.000 ;
    END
  END data_write_data[0]
  PIN data_write_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1342.880 996.000 1343.440 1000.000 ;
    END
  END data_write_data[10]
  PIN data_write_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1355.200 996.000 1355.760 1000.000 ;
    END
  END data_write_data[11]
  PIN data_write_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1367.520 996.000 1368.080 1000.000 ;
    END
  END data_write_data[12]
  PIN data_write_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1379.840 996.000 1380.400 1000.000 ;
    END
  END data_write_data[13]
  PIN data_write_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1392.160 996.000 1392.720 1000.000 ;
    END
  END data_write_data[14]
  PIN data_write_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1404.480 996.000 1405.040 1000.000 ;
    END
  END data_write_data[15]
  PIN data_write_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1151.920 996.000 1152.480 1000.000 ;
    END
  END data_write_data[1]
  PIN data_write_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1176.560 996.000 1177.120 1000.000 ;
    END
  END data_write_data[2]
  PIN data_write_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1201.200 996.000 1201.760 1000.000 ;
    END
  END data_write_data[3]
  PIN data_write_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1225.840 996.000 1226.400 1000.000 ;
    END
  END data_write_data[4]
  PIN data_write_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1250.480 996.000 1251.040 1000.000 ;
    END
  END data_write_data[5]
  PIN data_write_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1275.120 996.000 1275.680 1000.000 ;
    END
  END data_write_data[6]
  PIN data_write_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1299.760 996.000 1300.320 1000.000 ;
    END
  END data_write_data[7]
  PIN data_write_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1318.240 996.000 1318.800 1000.000 ;
    END
  END data_write_data[8]
  PIN data_write_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1330.560 996.000 1331.120 1000.000 ;
    END
  END data_write_data[9]
  PIN dataw_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1108.800 996.000 1109.360 1000.000 ;
    END
  END dataw_en
  PIN dataw_en_8bit[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1133.440 996.000 1134.000 1000.000 ;
    END
  END dataw_en_8bit[0]
  PIN dataw_en_8bit[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1158.080 996.000 1158.640 1000.000 ;
    END
  END dataw_en_8bit[1]
  PIN dataw_en_8bit[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1182.720 996.000 1183.280 1000.000 ;
    END
  END dataw_en_8bit[2]
  PIN dataw_en_8bit[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1207.360 996.000 1207.920 1000.000 ;
    END
  END dataw_en_8bit[3]
  PIN dataw_en_8bit[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1232.000 996.000 1232.560 1000.000 ;
    END
  END dataw_en_8bit[4]
  PIN dataw_en_8bit[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1256.640 996.000 1257.200 1000.000 ;
    END
  END dataw_en_8bit[5]
  PIN dataw_en_8bit[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1281.280 996.000 1281.840 1000.000 ;
    END
  END dataw_en_8bit[6]
  PIN dataw_en_8bit[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1305.920 996.000 1306.480 1000.000 ;
    END
  END dataw_en_8bit[7]
  PIN hlt
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1718.640 996.000 1719.200 1000.000 ;
    END
  END hlt
  PIN instr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1422.960 996.000 1423.520 1000.000 ;
    END
  END instr[0]
  PIN instr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1644.720 996.000 1645.280 1000.000 ;
    END
  END instr[10]
  PIN instr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1657.040 996.000 1657.600 1000.000 ;
    END
  END instr[11]
  PIN instr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1669.360 996.000 1669.920 1000.000 ;
    END
  END instr[12]
  PIN instr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1681.680 996.000 1682.240 1000.000 ;
    END
  END instr[13]
  PIN instr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1694.000 996.000 1694.560 1000.000 ;
    END
  END instr[14]
  PIN instr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1706.320 996.000 1706.880 1000.000 ;
    END
  END instr[15]
  PIN instr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1447.600 996.000 1448.160 1000.000 ;
    END
  END instr[1]
  PIN instr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1472.240 996.000 1472.800 1000.000 ;
    END
  END instr[2]
  PIN instr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1496.880 996.000 1497.440 1000.000 ;
    END
  END instr[3]
  PIN instr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1521.520 996.000 1522.080 1000.000 ;
    END
  END instr[4]
  PIN instr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1546.160 996.000 1546.720 1000.000 ;
    END
  END instr[5]
  PIN instr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1570.800 996.000 1571.360 1000.000 ;
    END
  END instr[6]
  PIN instr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1595.440 996.000 1596.000 1000.000 ;
    END
  END instr[7]
  PIN instr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1620.080 996.000 1620.640 1000.000 ;
    END
  END instr[8]
  PIN instr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1632.400 996.000 1632.960 1000.000 ;
    END
  END instr[9]
  PIN instr_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1429.120 996.000 1429.680 1000.000 ;
    END
  END instr_mem_addr[0]
  PIN instr_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1453.760 996.000 1454.320 1000.000 ;
    END
  END instr_mem_addr[1]
  PIN instr_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1478.400 996.000 1478.960 1000.000 ;
    END
  END instr_mem_addr[2]
  PIN instr_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1503.040 996.000 1503.600 1000.000 ;
    END
  END instr_mem_addr[3]
  PIN instr_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1527.680 996.000 1528.240 1000.000 ;
    END
  END instr_mem_addr[4]
  PIN instr_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1552.320 996.000 1552.880 1000.000 ;
    END
  END instr_mem_addr[5]
  PIN instr_mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1576.960 996.000 1577.520 1000.000 ;
    END
  END instr_mem_addr[6]
  PIN instr_mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1601.600 996.000 1602.160 1000.000 ;
    END
  END instr_mem_addr[7]
  PIN instr_mem_sel
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1410.640 996.000 1411.200 1000.000 ;
    END
  END instr_mem_sel
  PIN instr_write_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1435.280 996.000 1435.840 1000.000 ;
    END
  END instr_write_data[0]
  PIN instr_write_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1650.880 996.000 1651.440 1000.000 ;
    END
  END instr_write_data[10]
  PIN instr_write_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1663.200 996.000 1663.760 1000.000 ;
    END
  END instr_write_data[11]
  PIN instr_write_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1675.520 996.000 1676.080 1000.000 ;
    END
  END instr_write_data[12]
  PIN instr_write_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1687.840 996.000 1688.400 1000.000 ;
    END
  END instr_write_data[13]
  PIN instr_write_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1700.160 996.000 1700.720 1000.000 ;
    END
  END instr_write_data[14]
  PIN instr_write_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1712.480 996.000 1713.040 1000.000 ;
    END
  END instr_write_data[15]
  PIN instr_write_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1459.920 996.000 1460.480 1000.000 ;
    END
  END instr_write_data[1]
  PIN instr_write_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1484.560 996.000 1485.120 1000.000 ;
    END
  END instr_write_data[2]
  PIN instr_write_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1509.200 996.000 1509.760 1000.000 ;
    END
  END instr_write_data[3]
  PIN instr_write_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1533.840 996.000 1534.400 1000.000 ;
    END
  END instr_write_data[4]
  PIN instr_write_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1558.480 996.000 1559.040 1000.000 ;
    END
  END instr_write_data[5]
  PIN instr_write_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1583.120 996.000 1583.680 1000.000 ;
    END
  END instr_write_data[6]
  PIN instr_write_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1607.760 996.000 1608.320 1000.000 ;
    END
  END instr_write_data[7]
  PIN instr_write_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1626.240 996.000 1626.800 1000.000 ;
    END
  END instr_write_data[8]
  PIN instr_write_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1638.560 996.000 1639.120 1000.000 ;
    END
  END instr_write_data[9]
  PIN instrw_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1416.800 996.000 1417.360 1000.000 ;
    END
  END instrw_en
  PIN instrw_en_8bit[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1441.440 996.000 1442.000 1000.000 ;
    END
  END instrw_en_8bit[0]
  PIN instrw_en_8bit[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1466.080 996.000 1466.640 1000.000 ;
    END
  END instrw_en_8bit[1]
  PIN instrw_en_8bit[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1490.720 996.000 1491.280 1000.000 ;
    END
  END instrw_en_8bit[2]
  PIN instrw_en_8bit[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1515.360 996.000 1515.920 1000.000 ;
    END
  END instrw_en_8bit[3]
  PIN instrw_en_8bit[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1540.000 996.000 1540.560 1000.000 ;
    END
  END instrw_en_8bit[4]
  PIN instrw_en_8bit[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1564.640 996.000 1565.200 1000.000 ;
    END
  END instrw_en_8bit[5]
  PIN instrw_en_8bit[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1589.280 996.000 1589.840 1000.000 ;
    END
  END instrw_en_8bit[6]
  PIN instrw_en_8bit[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1613.920 996.000 1614.480 1000.000 ;
    END
  END instrw_en_8bit[7]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.760 996.000 68.320 1000.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 252.560 996.000 253.120 1000.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 271.040 996.000 271.600 1000.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 289.520 996.000 290.080 1000.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 308.000 996.000 308.560 1000.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 326.480 996.000 327.040 1000.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 344.960 996.000 345.520 1000.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 363.440 996.000 364.000 1000.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 381.920 996.000 382.480 1000.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 400.400 996.000 400.960 1000.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 418.880 996.000 419.440 1000.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 996.000 86.800 1000.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 437.360 996.000 437.920 1000.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 455.840 996.000 456.400 1000.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 474.320 996.000 474.880 1000.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 492.800 996.000 493.360 1000.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 511.280 996.000 511.840 1000.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 529.760 996.000 530.320 1000.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 548.240 996.000 548.800 1000.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 566.720 996.000 567.280 1000.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 585.200 996.000 585.760 1000.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 603.680 996.000 604.240 1000.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.720 996.000 105.280 1000.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 622.160 996.000 622.720 1000.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 640.640 996.000 641.200 1000.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 659.120 996.000 659.680 1000.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 677.600 996.000 678.160 1000.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 696.080 996.000 696.640 1000.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 714.560 996.000 715.120 1000.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 733.040 996.000 733.600 1000.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 751.520 996.000 752.080 1000.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 996.000 123.760 1000.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 141.680 996.000 142.240 1000.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 160.160 996.000 160.720 1000.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 178.640 996.000 179.200 1000.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 197.120 996.000 197.680 1000.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.600 996.000 216.160 1000.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.080 996.000 234.640 1000.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 996.000 74.480 1000.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 996.000 259.280 1000.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 277.200 996.000 277.760 1000.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 295.680 996.000 296.240 1000.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 314.160 996.000 314.720 1000.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 332.640 996.000 333.200 1000.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 351.120 996.000 351.680 1000.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 369.600 996.000 370.160 1000.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 388.080 996.000 388.640 1000.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 996.000 407.120 1000.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 425.040 996.000 425.600 1000.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 92.400 996.000 92.960 1000.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 443.520 996.000 444.080 1000.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 462.000 996.000 462.560 1000.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 480.480 996.000 481.040 1000.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 498.960 996.000 499.520 1000.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 996.000 518.000 1000.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 535.920 996.000 536.480 1000.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 554.400 996.000 554.960 1000.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 572.880 996.000 573.440 1000.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 591.360 996.000 591.920 1000.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 609.840 996.000 610.400 1000.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 996.000 111.440 1000.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 628.320 996.000 628.880 1000.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 646.800 996.000 647.360 1000.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 665.280 996.000 665.840 1000.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 683.760 996.000 684.320 1000.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 702.240 996.000 702.800 1000.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 720.720 996.000 721.280 1000.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 739.200 996.000 739.760 1000.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 757.680 996.000 758.240 1000.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 129.360 996.000 129.920 1000.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 996.000 148.400 1000.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 166.320 996.000 166.880 1000.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 996.000 185.360 1000.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 203.280 996.000 203.840 1000.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 996.000 222.320 1000.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 240.240 996.000 240.800 1000.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 80.080 996.000 80.640 1000.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 264.880 996.000 265.440 1000.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 283.360 996.000 283.920 1000.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 301.840 996.000 302.400 1000.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 320.320 996.000 320.880 1000.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 338.800 996.000 339.360 1000.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 357.280 996.000 357.840 1000.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 375.760 996.000 376.320 1000.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 394.240 996.000 394.800 1000.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 412.720 996.000 413.280 1000.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 431.200 996.000 431.760 1000.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 996.000 99.120 1000.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 449.680 996.000 450.240 1000.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 468.160 996.000 468.720 1000.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 486.640 996.000 487.200 1000.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 505.120 996.000 505.680 1000.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 523.600 996.000 524.160 1000.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 542.080 996.000 542.640 1000.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 560.560 996.000 561.120 1000.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 579.040 996.000 579.600 1000.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 597.520 996.000 598.080 1000.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 616.000 996.000 616.560 1000.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.040 996.000 117.600 1000.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 634.480 996.000 635.040 1000.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 652.960 996.000 653.520 1000.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 671.440 996.000 672.000 1000.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 689.920 996.000 690.480 1000.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 708.400 996.000 708.960 1000.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 726.880 996.000 727.440 1000.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 745.360 996.000 745.920 1000.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 763.840 996.000 764.400 1000.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 996.000 136.080 1000.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.000 996.000 154.560 1000.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 172.480 996.000 173.040 1000.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 190.960 996.000 191.520 1000.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 209.440 996.000 210.000 1000.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 227.920 996.000 228.480 1000.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 246.400 996.000 246.960 1000.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1762.880 0.000 1763.440 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1766.240 0.000 1766.800 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1769.600 0.000 1770.160 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 375.200 0.000 375.760 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1383.200 0.000 1383.760 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1393.280 0.000 1393.840 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1403.360 0.000 1403.920 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1413.440 0.000 1414.000 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1423.520 0.000 1424.080 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1433.600 0.000 1434.160 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1443.680 0.000 1444.240 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1453.760 0.000 1454.320 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1463.840 0.000 1464.400 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1473.920 0.000 1474.480 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 476.000 0.000 476.560 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1484.000 0.000 1484.560 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1494.080 0.000 1494.640 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1504.160 0.000 1504.720 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1514.240 0.000 1514.800 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1524.320 0.000 1524.880 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1534.400 0.000 1534.960 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1544.480 0.000 1545.040 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1554.560 0.000 1555.120 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1564.640 0.000 1565.200 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1574.720 0.000 1575.280 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 486.080 0.000 486.640 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1584.800 0.000 1585.360 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1594.880 0.000 1595.440 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1604.960 0.000 1605.520 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1615.040 0.000 1615.600 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1625.120 0.000 1625.680 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1635.200 0.000 1635.760 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1645.280 0.000 1645.840 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1655.360 0.000 1655.920 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 496.160 0.000 496.720 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 506.240 0.000 506.800 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 516.320 0.000 516.880 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 526.400 0.000 526.960 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 536.480 0.000 537.040 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 546.560 0.000 547.120 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 556.640 0.000 557.200 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 566.720 0.000 567.280 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 385.280 0.000 385.840 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 576.800 0.000 577.360 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 586.880 0.000 587.440 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 596.960 0.000 597.520 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 607.040 0.000 607.600 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 617.120 0.000 617.680 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 627.200 0.000 627.760 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 637.280 0.000 637.840 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 647.360 0.000 647.920 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 657.440 0.000 658.000 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 667.520 0.000 668.080 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 395.360 0.000 395.920 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 677.600 0.000 678.160 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 687.680 0.000 688.240 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 697.760 0.000 698.320 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 707.840 0.000 708.400 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 717.920 0.000 718.480 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 728.000 0.000 728.560 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 738.080 0.000 738.640 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 748.160 0.000 748.720 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 758.240 0.000 758.800 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 768.320 0.000 768.880 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 405.440 0.000 406.000 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 778.400 0.000 778.960 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 788.480 0.000 789.040 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 798.560 0.000 799.120 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 808.640 0.000 809.200 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 818.720 0.000 819.280 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 828.800 0.000 829.360 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 838.880 0.000 839.440 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 848.960 0.000 849.520 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 859.040 0.000 859.600 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 869.120 0.000 869.680 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 415.520 0.000 416.080 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 879.200 0.000 879.760 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 889.280 0.000 889.840 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 899.360 0.000 899.920 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 909.440 0.000 910.000 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 919.520 0.000 920.080 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 929.600 0.000 930.160 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 939.680 0.000 940.240 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 949.760 0.000 950.320 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 959.840 0.000 960.400 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 969.920 0.000 970.480 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 425.600 0.000 426.160 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 980.000 0.000 980.560 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 990.080 0.000 990.640 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1000.160 0.000 1000.720 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1010.240 0.000 1010.800 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1020.320 0.000 1020.880 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1030.400 0.000 1030.960 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1040.480 0.000 1041.040 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1050.560 0.000 1051.120 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1060.640 0.000 1061.200 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1070.720 0.000 1071.280 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 435.680 0.000 436.240 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1080.800 0.000 1081.360 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1090.880 0.000 1091.440 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1100.960 0.000 1101.520 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1111.040 0.000 1111.600 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1121.120 0.000 1121.680 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1131.200 0.000 1131.760 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1141.280 0.000 1141.840 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1151.360 0.000 1151.920 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1161.440 0.000 1162.000 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1171.520 0.000 1172.080 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 445.760 0.000 446.320 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1181.600 0.000 1182.160 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1191.680 0.000 1192.240 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1201.760 0.000 1202.320 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1211.840 0.000 1212.400 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1221.920 0.000 1222.480 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1232.000 0.000 1232.560 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1242.080 0.000 1242.640 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1252.160 0.000 1252.720 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1262.240 0.000 1262.800 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1272.320 0.000 1272.880 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 455.840 0.000 456.400 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1282.400 0.000 1282.960 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1292.480 0.000 1293.040 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1302.560 0.000 1303.120 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1312.640 0.000 1313.200 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1322.720 0.000 1323.280 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1332.800 0.000 1333.360 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1342.880 0.000 1343.440 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1352.960 0.000 1353.520 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1363.040 0.000 1363.600 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1373.120 0.000 1373.680 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 465.920 0.000 466.480 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 378.560 0.000 379.120 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1386.560 0.000 1387.120 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1396.640 0.000 1397.200 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1406.720 0.000 1407.280 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1416.800 0.000 1417.360 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1426.880 0.000 1427.440 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1436.960 0.000 1437.520 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1447.040 0.000 1447.600 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1457.120 0.000 1457.680 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1467.200 0.000 1467.760 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1477.280 0.000 1477.840 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 479.360 0.000 479.920 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1487.360 0.000 1487.920 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1497.440 0.000 1498.000 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1507.520 0.000 1508.080 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1517.600 0.000 1518.160 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1527.680 0.000 1528.240 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1537.760 0.000 1538.320 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1547.840 0.000 1548.400 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1557.920 0.000 1558.480 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1568.000 0.000 1568.560 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1578.080 0.000 1578.640 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 489.440 0.000 490.000 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1588.160 0.000 1588.720 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1598.240 0.000 1598.800 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1608.320 0.000 1608.880 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1618.400 0.000 1618.960 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1628.480 0.000 1629.040 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1638.560 0.000 1639.120 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1648.640 0.000 1649.200 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1658.720 0.000 1659.280 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 499.520 0.000 500.080 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 509.600 0.000 510.160 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 519.680 0.000 520.240 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 529.760 0.000 530.320 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 539.840 0.000 540.400 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 549.920 0.000 550.480 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 560.000 0.000 560.560 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 570.080 0.000 570.640 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 388.640 0.000 389.200 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 580.160 0.000 580.720 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 590.240 0.000 590.800 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 600.320 0.000 600.880 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 610.400 0.000 610.960 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 620.480 0.000 621.040 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 630.560 0.000 631.120 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 640.640 0.000 641.200 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 650.720 0.000 651.280 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 660.800 0.000 661.360 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 670.880 0.000 671.440 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 398.720 0.000 399.280 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 680.960 0.000 681.520 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 691.040 0.000 691.600 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 701.120 0.000 701.680 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 711.200 0.000 711.760 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 721.280 0.000 721.840 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 731.360 0.000 731.920 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 741.440 0.000 742.000 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 751.520 0.000 752.080 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 761.600 0.000 762.160 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 771.680 0.000 772.240 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 408.800 0.000 409.360 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 781.760 0.000 782.320 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 791.840 0.000 792.400 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 801.920 0.000 802.480 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 812.000 0.000 812.560 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 822.080 0.000 822.640 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 832.160 0.000 832.720 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 842.240 0.000 842.800 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 852.320 0.000 852.880 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 862.400 0.000 862.960 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 872.480 0.000 873.040 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 418.880 0.000 419.440 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 882.560 0.000 883.120 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 892.640 0.000 893.200 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 902.720 0.000 903.280 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 912.800 0.000 913.360 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 922.880 0.000 923.440 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 932.960 0.000 933.520 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 943.040 0.000 943.600 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 953.120 0.000 953.680 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 963.200 0.000 963.760 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 973.280 0.000 973.840 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 428.960 0.000 429.520 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 983.360 0.000 983.920 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 993.440 0.000 994.000 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1003.520 0.000 1004.080 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1013.600 0.000 1014.160 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1023.680 0.000 1024.240 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1033.760 0.000 1034.320 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1043.840 0.000 1044.400 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1053.920 0.000 1054.480 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1064.000 0.000 1064.560 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1074.080 0.000 1074.640 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 439.040 0.000 439.600 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1084.160 0.000 1084.720 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1094.240 0.000 1094.800 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1104.320 0.000 1104.880 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1114.400 0.000 1114.960 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1124.480 0.000 1125.040 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1134.560 0.000 1135.120 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1144.640 0.000 1145.200 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1154.720 0.000 1155.280 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1164.800 0.000 1165.360 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1174.880 0.000 1175.440 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 449.120 0.000 449.680 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1184.960 0.000 1185.520 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1195.040 0.000 1195.600 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1205.120 0.000 1205.680 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1215.200 0.000 1215.760 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1225.280 0.000 1225.840 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1235.360 0.000 1235.920 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1245.440 0.000 1246.000 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1255.520 0.000 1256.080 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1265.600 0.000 1266.160 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1275.680 0.000 1276.240 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 459.200 0.000 459.760 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1285.760 0.000 1286.320 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1295.840 0.000 1296.400 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1305.920 0.000 1306.480 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1316.000 0.000 1316.560 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1326.080 0.000 1326.640 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1336.160 0.000 1336.720 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1346.240 0.000 1346.800 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1356.320 0.000 1356.880 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1366.400 0.000 1366.960 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1376.480 0.000 1377.040 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 469.280 0.000 469.840 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 381.920 0.000 382.480 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1389.920 0.000 1390.480 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1400.000 0.000 1400.560 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1410.080 0.000 1410.640 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1420.160 0.000 1420.720 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1430.240 0.000 1430.800 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1440.320 0.000 1440.880 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1450.400 0.000 1450.960 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1460.480 0.000 1461.040 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1470.560 0.000 1471.120 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1480.640 0.000 1481.200 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 482.720 0.000 483.280 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1490.720 0.000 1491.280 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1500.800 0.000 1501.360 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1510.880 0.000 1511.440 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1520.960 0.000 1521.520 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1531.040 0.000 1531.600 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1541.120 0.000 1541.680 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1551.200 0.000 1551.760 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1561.280 0.000 1561.840 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1571.360 0.000 1571.920 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1581.440 0.000 1582.000 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 492.800 0.000 493.360 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1591.520 0.000 1592.080 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1601.600 0.000 1602.160 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1611.680 0.000 1612.240 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1621.760 0.000 1622.320 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1631.840 0.000 1632.400 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1641.920 0.000 1642.480 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1652.000 0.000 1652.560 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1662.080 0.000 1662.640 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 502.880 0.000 503.440 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 512.960 0.000 513.520 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 523.040 0.000 523.600 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 533.120 0.000 533.680 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 543.200 0.000 543.760 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 553.280 0.000 553.840 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 563.360 0.000 563.920 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 573.440 0.000 574.000 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 392.000 0.000 392.560 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 583.520 0.000 584.080 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 593.600 0.000 594.160 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 603.680 0.000 604.240 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 613.760 0.000 614.320 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 623.840 0.000 624.400 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 633.920 0.000 634.480 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 644.000 0.000 644.560 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 654.080 0.000 654.640 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 664.160 0.000 664.720 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 674.240 0.000 674.800 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 402.080 0.000 402.640 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 684.320 0.000 684.880 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 694.400 0.000 694.960 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 704.480 0.000 705.040 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 714.560 0.000 715.120 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 724.640 0.000 725.200 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 734.720 0.000 735.280 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 744.800 0.000 745.360 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 754.880 0.000 755.440 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 764.960 0.000 765.520 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 775.040 0.000 775.600 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 412.160 0.000 412.720 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 785.120 0.000 785.680 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 795.200 0.000 795.760 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 805.280 0.000 805.840 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 815.360 0.000 815.920 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 825.440 0.000 826.000 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 835.520 0.000 836.080 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 845.600 0.000 846.160 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 855.680 0.000 856.240 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 865.760 0.000 866.320 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 875.840 0.000 876.400 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 422.240 0.000 422.800 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 885.920 0.000 886.480 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 896.000 0.000 896.560 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 906.080 0.000 906.640 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 916.160 0.000 916.720 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 926.240 0.000 926.800 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 936.320 0.000 936.880 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 946.400 0.000 946.960 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 956.480 0.000 957.040 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 966.560 0.000 967.120 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 976.640 0.000 977.200 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 432.320 0.000 432.880 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 986.720 0.000 987.280 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 996.800 0.000 997.360 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1006.880 0.000 1007.440 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1016.960 0.000 1017.520 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1027.040 0.000 1027.600 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1037.120 0.000 1037.680 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1047.200 0.000 1047.760 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1057.280 0.000 1057.840 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1067.360 0.000 1067.920 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1077.440 0.000 1078.000 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 442.400 0.000 442.960 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1087.520 0.000 1088.080 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1097.600 0.000 1098.160 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1107.680 0.000 1108.240 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1117.760 0.000 1118.320 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1127.840 0.000 1128.400 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1137.920 0.000 1138.480 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1148.000 0.000 1148.560 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1158.080 0.000 1158.640 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1168.160 0.000 1168.720 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1178.240 0.000 1178.800 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 452.480 0.000 453.040 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1188.320 0.000 1188.880 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1198.400 0.000 1198.960 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1208.480 0.000 1209.040 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1218.560 0.000 1219.120 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1228.640 0.000 1229.200 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1238.720 0.000 1239.280 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1248.800 0.000 1249.360 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1258.880 0.000 1259.440 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1268.960 0.000 1269.520 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1279.040 0.000 1279.600 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 462.560 0.000 463.120 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1289.120 0.000 1289.680 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1299.200 0.000 1299.760 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1309.280 0.000 1309.840 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1319.360 0.000 1319.920 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1329.440 0.000 1330.000 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1339.520 0.000 1340.080 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1349.600 0.000 1350.160 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1359.680 0.000 1360.240 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1369.760 0.000 1370.320 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1379.840 0.000 1380.400 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 472.640 0.000 473.200 4.000 ;
    END
  END la_oenb[9]
  PIN reset
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1779.680 0.000 1780.240 4.000 ;
    END
  END reset
  PIN start
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1776.320 0.000 1776.880 4.000 ;
    END
  END start
  PIN uP_data_mem_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 776.160 996.000 776.720 1000.000 ;
    END
  END uP_data_mem_addr[0]
  PIN uP_data_mem_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 800.800 996.000 801.360 1000.000 ;
    END
  END uP_data_mem_addr[1]
  PIN uP_data_mem_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 825.440 996.000 826.000 1000.000 ;
    END
  END uP_data_mem_addr[2]
  PIN uP_data_mem_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 850.080 996.000 850.640 1000.000 ;
    END
  END uP_data_mem_addr[3]
  PIN uP_data_mem_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 874.720 996.000 875.280 1000.000 ;
    END
  END uP_data_mem_addr[4]
  PIN uP_data_mem_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 899.360 996.000 899.920 1000.000 ;
    END
  END uP_data_mem_addr[5]
  PIN uP_data_mem_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 924.000 996.000 924.560 1000.000 ;
    END
  END uP_data_mem_addr[6]
  PIN uP_data_mem_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 948.640 996.000 949.200 1000.000 ;
    END
  END uP_data_mem_addr[7]
  PIN uP_dataw_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 770.000 996.000 770.560 1000.000 ;
    END
  END uP_dataw_en
  PIN uP_instr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 782.320 996.000 782.880 1000.000 ;
    END
  END uP_instr[0]
  PIN uP_instr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1010.240 996.000 1010.800 1000.000 ;
    END
  END uP_instr[10]
  PIN uP_instr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1028.720 996.000 1029.280 1000.000 ;
    END
  END uP_instr[11]
  PIN uP_instr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1047.200 996.000 1047.760 1000.000 ;
    END
  END uP_instr[12]
  PIN uP_instr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1065.680 996.000 1066.240 1000.000 ;
    END
  END uP_instr[13]
  PIN uP_instr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1078.000 996.000 1078.560 1000.000 ;
    END
  END uP_instr[14]
  PIN uP_instr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1090.320 996.000 1090.880 1000.000 ;
    END
  END uP_instr[15]
  PIN uP_instr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 806.960 996.000 807.520 1000.000 ;
    END
  END uP_instr[1]
  PIN uP_instr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 831.600 996.000 832.160 1000.000 ;
    END
  END uP_instr[2]
  PIN uP_instr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 856.240 996.000 856.800 1000.000 ;
    END
  END uP_instr[3]
  PIN uP_instr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 880.880 996.000 881.440 1000.000 ;
    END
  END uP_instr[4]
  PIN uP_instr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 905.520 996.000 906.080 1000.000 ;
    END
  END uP_instr[5]
  PIN uP_instr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 930.160 996.000 930.720 1000.000 ;
    END
  END uP_instr[6]
  PIN uP_instr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 954.800 996.000 955.360 1000.000 ;
    END
  END uP_instr[7]
  PIN uP_instr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 973.280 996.000 973.840 1000.000 ;
    END
  END uP_instr[8]
  PIN uP_instr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 991.760 996.000 992.320 1000.000 ;
    END
  END uP_instr[9]
  PIN uP_instr_mem_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 788.480 996.000 789.040 1000.000 ;
    END
  END uP_instr_mem_addr[0]
  PIN uP_instr_mem_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1016.400 996.000 1016.960 1000.000 ;
    END
  END uP_instr_mem_addr[10]
  PIN uP_instr_mem_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1034.880 996.000 1035.440 1000.000 ;
    END
  END uP_instr_mem_addr[11]
  PIN uP_instr_mem_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1053.360 996.000 1053.920 1000.000 ;
    END
  END uP_instr_mem_addr[12]
  PIN uP_instr_mem_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 813.120 996.000 813.680 1000.000 ;
    END
  END uP_instr_mem_addr[1]
  PIN uP_instr_mem_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 837.760 996.000 838.320 1000.000 ;
    END
  END uP_instr_mem_addr[2]
  PIN uP_instr_mem_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 862.400 996.000 862.960 1000.000 ;
    END
  END uP_instr_mem_addr[3]
  PIN uP_instr_mem_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 887.040 996.000 887.600 1000.000 ;
    END
  END uP_instr_mem_addr[4]
  PIN uP_instr_mem_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 911.680 996.000 912.240 1000.000 ;
    END
  END uP_instr_mem_addr[5]
  PIN uP_instr_mem_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 936.320 996.000 936.880 1000.000 ;
    END
  END uP_instr_mem_addr[6]
  PIN uP_instr_mem_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 960.960 996.000 961.520 1000.000 ;
    END
  END uP_instr_mem_addr[7]
  PIN uP_instr_mem_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 979.440 996.000 980.000 1000.000 ;
    END
  END uP_instr_mem_addr[8]
  PIN uP_instr_mem_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 997.920 996.000 998.480 1000.000 ;
    END
  END uP_instr_mem_addr[9]
  PIN uP_write_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 794.640 996.000 795.200 1000.000 ;
    END
  END uP_write_data[0]
  PIN uP_write_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1022.560 996.000 1023.120 1000.000 ;
    END
  END uP_write_data[10]
  PIN uP_write_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1041.040 996.000 1041.600 1000.000 ;
    END
  END uP_write_data[11]
  PIN uP_write_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1059.520 996.000 1060.080 1000.000 ;
    END
  END uP_write_data[12]
  PIN uP_write_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1071.840 996.000 1072.400 1000.000 ;
    END
  END uP_write_data[13]
  PIN uP_write_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1084.160 996.000 1084.720 1000.000 ;
    END
  END uP_write_data[14]
  PIN uP_write_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1096.480 996.000 1097.040 1000.000 ;
    END
  END uP_write_data[15]
  PIN uP_write_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 819.280 996.000 819.840 1000.000 ;
    END
  END uP_write_data[1]
  PIN uP_write_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 843.920 996.000 844.480 1000.000 ;
    END
  END uP_write_data[2]
  PIN uP_write_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 868.560 996.000 869.120 1000.000 ;
    END
  END uP_write_data[3]
  PIN uP_write_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 893.200 996.000 893.760 1000.000 ;
    END
  END uP_write_data[4]
  PIN uP_write_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 917.840 996.000 918.400 1000.000 ;
    END
  END uP_write_data[5]
  PIN uP_write_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 942.480 996.000 943.040 1000.000 ;
    END
  END uP_write_data[6]
  PIN uP_write_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 967.120 996.000 967.680 1000.000 ;
    END
  END uP_write_data[7]
  PIN uP_write_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 985.600 996.000 986.160 1000.000 ;
    END
  END uP_write_data[8]
  PIN uP_write_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1004.080 996.000 1004.640 1000.000 ;
    END
  END uP_write_data[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1558.240 15.380 1559.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1711.840 15.380 1713.440 984.220 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.040 15.380 1636.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.640 15.380 1790.240 984.220 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 19.040 0.000 19.600 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 22.400 0.000 22.960 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 25.760 0.000 26.320 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 39.200 0.000 39.760 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 153.440 0.000 154.000 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 163.520 0.000 164.080 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 173.600 0.000 174.160 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 183.680 0.000 184.240 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 193.760 0.000 194.320 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 203.840 0.000 204.400 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 213.920 0.000 214.480 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 224.000 0.000 224.560 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 234.080 0.000 234.640 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 244.160 0.000 244.720 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 52.640 0.000 53.200 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 254.240 0.000 254.800 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 264.320 0.000 264.880 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 274.400 0.000 274.960 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 284.480 0.000 285.040 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 294.560 0.000 295.120 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 304.640 0.000 305.200 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 314.720 0.000 315.280 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 324.800 0.000 325.360 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 334.880 0.000 335.440 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 344.960 0.000 345.520 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 0.000 66.640 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 355.040 0.000 355.600 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 365.120 0.000 365.680 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 79.520 0.000 80.080 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 92.960 0.000 93.520 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 103.040 0.000 103.600 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 0.000 113.680 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 123.200 0.000 123.760 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 133.280 0.000 133.840 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 143.360 0.000 143.920 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.120 0.000 29.680 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 42.560 0.000 43.120 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 156.800 0.000 157.360 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 0.000 167.440 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 176.960 0.000 177.520 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 187.040 0.000 187.600 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 197.120 0.000 197.680 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 207.200 0.000 207.760 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 217.280 0.000 217.840 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 227.360 0.000 227.920 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 237.440 0.000 238.000 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 247.520 0.000 248.080 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 56.000 0.000 56.560 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 257.600 0.000 258.160 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 267.680 0.000 268.240 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 277.760 0.000 278.320 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 287.840 0.000 288.400 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 297.920 0.000 298.480 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 308.000 0.000 308.560 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 318.080 0.000 318.640 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 328.160 0.000 328.720 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 338.240 0.000 338.800 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 348.320 0.000 348.880 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 69.440 0.000 70.000 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 358.400 0.000 358.960 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 368.480 0.000 369.040 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 82.880 0.000 83.440 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 0.000 96.880 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 0.000 106.960 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 0.000 117.040 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 0.000 127.120 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 136.640 0.000 137.200 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 0.000 147.280 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 0.000 46.480 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 160.160 0.000 160.720 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 170.240 0.000 170.800 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 180.320 0.000 180.880 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 190.400 0.000 190.960 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 200.480 0.000 201.040 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 210.560 0.000 211.120 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 220.640 0.000 221.200 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 230.720 0.000 231.280 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 240.800 0.000 241.360 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 250.880 0.000 251.440 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 0.000 59.920 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 260.960 0.000 261.520 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 271.040 0.000 271.600 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.120 0.000 281.680 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 291.200 0.000 291.760 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 301.280 0.000 301.840 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 311.360 0.000 311.920 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 321.440 0.000 322.000 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 331.520 0.000 332.080 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 341.600 0.000 342.160 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 351.680 0.000 352.240 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 72.800 0.000 73.360 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 361.760 0.000 362.320 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 371.840 0.000 372.400 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 0.000 86.800 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 99.680 0.000 100.240 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 109.760 0.000 110.320 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 119.840 0.000 120.400 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 129.920 0.000 130.480 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 0.000 140.560 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 150.080 0.000 150.640 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 49.280 0.000 49.840 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 62.720 0.000 63.280 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 76.160 0.000 76.720 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 89.600 0.000 90.160 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 32.480 0.000 33.040 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 35.840 0.000 36.400 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 14.150 1793.120 984.890 ;
      LAYER Metal2 ;
        RECT 16.380 995.700 67.460 997.830 ;
        RECT 68.620 995.700 73.620 997.830 ;
        RECT 74.780 995.700 79.780 997.830 ;
        RECT 80.940 995.700 85.940 997.830 ;
        RECT 87.100 995.700 92.100 997.830 ;
        RECT 93.260 995.700 98.260 997.830 ;
        RECT 99.420 995.700 104.420 997.830 ;
        RECT 105.580 995.700 110.580 997.830 ;
        RECT 111.740 995.700 116.740 997.830 ;
        RECT 117.900 995.700 122.900 997.830 ;
        RECT 124.060 995.700 129.060 997.830 ;
        RECT 130.220 995.700 135.220 997.830 ;
        RECT 136.380 995.700 141.380 997.830 ;
        RECT 142.540 995.700 147.540 997.830 ;
        RECT 148.700 995.700 153.700 997.830 ;
        RECT 154.860 995.700 159.860 997.830 ;
        RECT 161.020 995.700 166.020 997.830 ;
        RECT 167.180 995.700 172.180 997.830 ;
        RECT 173.340 995.700 178.340 997.830 ;
        RECT 179.500 995.700 184.500 997.830 ;
        RECT 185.660 995.700 190.660 997.830 ;
        RECT 191.820 995.700 196.820 997.830 ;
        RECT 197.980 995.700 202.980 997.830 ;
        RECT 204.140 995.700 209.140 997.830 ;
        RECT 210.300 995.700 215.300 997.830 ;
        RECT 216.460 995.700 221.460 997.830 ;
        RECT 222.620 995.700 227.620 997.830 ;
        RECT 228.780 995.700 233.780 997.830 ;
        RECT 234.940 995.700 239.940 997.830 ;
        RECT 241.100 995.700 246.100 997.830 ;
        RECT 247.260 995.700 252.260 997.830 ;
        RECT 253.420 995.700 258.420 997.830 ;
        RECT 259.580 995.700 264.580 997.830 ;
        RECT 265.740 995.700 270.740 997.830 ;
        RECT 271.900 995.700 276.900 997.830 ;
        RECT 278.060 995.700 283.060 997.830 ;
        RECT 284.220 995.700 289.220 997.830 ;
        RECT 290.380 995.700 295.380 997.830 ;
        RECT 296.540 995.700 301.540 997.830 ;
        RECT 302.700 995.700 307.700 997.830 ;
        RECT 308.860 995.700 313.860 997.830 ;
        RECT 315.020 995.700 320.020 997.830 ;
        RECT 321.180 995.700 326.180 997.830 ;
        RECT 327.340 995.700 332.340 997.830 ;
        RECT 333.500 995.700 338.500 997.830 ;
        RECT 339.660 995.700 344.660 997.830 ;
        RECT 345.820 995.700 350.820 997.830 ;
        RECT 351.980 995.700 356.980 997.830 ;
        RECT 358.140 995.700 363.140 997.830 ;
        RECT 364.300 995.700 369.300 997.830 ;
        RECT 370.460 995.700 375.460 997.830 ;
        RECT 376.620 995.700 381.620 997.830 ;
        RECT 382.780 995.700 387.780 997.830 ;
        RECT 388.940 995.700 393.940 997.830 ;
        RECT 395.100 995.700 400.100 997.830 ;
        RECT 401.260 995.700 406.260 997.830 ;
        RECT 407.420 995.700 412.420 997.830 ;
        RECT 413.580 995.700 418.580 997.830 ;
        RECT 419.740 995.700 424.740 997.830 ;
        RECT 425.900 995.700 430.900 997.830 ;
        RECT 432.060 995.700 437.060 997.830 ;
        RECT 438.220 995.700 443.220 997.830 ;
        RECT 444.380 995.700 449.380 997.830 ;
        RECT 450.540 995.700 455.540 997.830 ;
        RECT 456.700 995.700 461.700 997.830 ;
        RECT 462.860 995.700 467.860 997.830 ;
        RECT 469.020 995.700 474.020 997.830 ;
        RECT 475.180 995.700 480.180 997.830 ;
        RECT 481.340 995.700 486.340 997.830 ;
        RECT 487.500 995.700 492.500 997.830 ;
        RECT 493.660 995.700 498.660 997.830 ;
        RECT 499.820 995.700 504.820 997.830 ;
        RECT 505.980 995.700 510.980 997.830 ;
        RECT 512.140 995.700 517.140 997.830 ;
        RECT 518.300 995.700 523.300 997.830 ;
        RECT 524.460 995.700 529.460 997.830 ;
        RECT 530.620 995.700 535.620 997.830 ;
        RECT 536.780 995.700 541.780 997.830 ;
        RECT 542.940 995.700 547.940 997.830 ;
        RECT 549.100 995.700 554.100 997.830 ;
        RECT 555.260 995.700 560.260 997.830 ;
        RECT 561.420 995.700 566.420 997.830 ;
        RECT 567.580 995.700 572.580 997.830 ;
        RECT 573.740 995.700 578.740 997.830 ;
        RECT 579.900 995.700 584.900 997.830 ;
        RECT 586.060 995.700 591.060 997.830 ;
        RECT 592.220 995.700 597.220 997.830 ;
        RECT 598.380 995.700 603.380 997.830 ;
        RECT 604.540 995.700 609.540 997.830 ;
        RECT 610.700 995.700 615.700 997.830 ;
        RECT 616.860 995.700 621.860 997.830 ;
        RECT 623.020 995.700 628.020 997.830 ;
        RECT 629.180 995.700 634.180 997.830 ;
        RECT 635.340 995.700 640.340 997.830 ;
        RECT 641.500 995.700 646.500 997.830 ;
        RECT 647.660 995.700 652.660 997.830 ;
        RECT 653.820 995.700 658.820 997.830 ;
        RECT 659.980 995.700 664.980 997.830 ;
        RECT 666.140 995.700 671.140 997.830 ;
        RECT 672.300 995.700 677.300 997.830 ;
        RECT 678.460 995.700 683.460 997.830 ;
        RECT 684.620 995.700 689.620 997.830 ;
        RECT 690.780 995.700 695.780 997.830 ;
        RECT 696.940 995.700 701.940 997.830 ;
        RECT 703.100 995.700 708.100 997.830 ;
        RECT 709.260 995.700 714.260 997.830 ;
        RECT 715.420 995.700 720.420 997.830 ;
        RECT 721.580 995.700 726.580 997.830 ;
        RECT 727.740 995.700 732.740 997.830 ;
        RECT 733.900 995.700 738.900 997.830 ;
        RECT 740.060 995.700 745.060 997.830 ;
        RECT 746.220 995.700 751.220 997.830 ;
        RECT 752.380 995.700 757.380 997.830 ;
        RECT 758.540 995.700 763.540 997.830 ;
        RECT 764.700 995.700 769.700 997.830 ;
        RECT 770.860 995.700 775.860 997.830 ;
        RECT 777.020 995.700 782.020 997.830 ;
        RECT 783.180 995.700 788.180 997.830 ;
        RECT 789.340 995.700 794.340 997.830 ;
        RECT 795.500 995.700 800.500 997.830 ;
        RECT 801.660 995.700 806.660 997.830 ;
        RECT 807.820 995.700 812.820 997.830 ;
        RECT 813.980 995.700 818.980 997.830 ;
        RECT 820.140 995.700 825.140 997.830 ;
        RECT 826.300 995.700 831.300 997.830 ;
        RECT 832.460 995.700 837.460 997.830 ;
        RECT 838.620 995.700 843.620 997.830 ;
        RECT 844.780 995.700 849.780 997.830 ;
        RECT 850.940 995.700 855.940 997.830 ;
        RECT 857.100 995.700 862.100 997.830 ;
        RECT 863.260 995.700 868.260 997.830 ;
        RECT 869.420 995.700 874.420 997.830 ;
        RECT 875.580 995.700 880.580 997.830 ;
        RECT 881.740 995.700 886.740 997.830 ;
        RECT 887.900 995.700 892.900 997.830 ;
        RECT 894.060 995.700 899.060 997.830 ;
        RECT 900.220 995.700 905.220 997.830 ;
        RECT 906.380 995.700 911.380 997.830 ;
        RECT 912.540 995.700 917.540 997.830 ;
        RECT 918.700 995.700 923.700 997.830 ;
        RECT 924.860 995.700 929.860 997.830 ;
        RECT 931.020 995.700 936.020 997.830 ;
        RECT 937.180 995.700 942.180 997.830 ;
        RECT 943.340 995.700 948.340 997.830 ;
        RECT 949.500 995.700 954.500 997.830 ;
        RECT 955.660 995.700 960.660 997.830 ;
        RECT 961.820 995.700 966.820 997.830 ;
        RECT 967.980 995.700 972.980 997.830 ;
        RECT 974.140 995.700 979.140 997.830 ;
        RECT 980.300 995.700 985.300 997.830 ;
        RECT 986.460 995.700 991.460 997.830 ;
        RECT 992.620 995.700 997.620 997.830 ;
        RECT 998.780 995.700 1003.780 997.830 ;
        RECT 1004.940 995.700 1009.940 997.830 ;
        RECT 1011.100 995.700 1016.100 997.830 ;
        RECT 1017.260 995.700 1022.260 997.830 ;
        RECT 1023.420 995.700 1028.420 997.830 ;
        RECT 1029.580 995.700 1034.580 997.830 ;
        RECT 1035.740 995.700 1040.740 997.830 ;
        RECT 1041.900 995.700 1046.900 997.830 ;
        RECT 1048.060 995.700 1053.060 997.830 ;
        RECT 1054.220 995.700 1059.220 997.830 ;
        RECT 1060.380 995.700 1065.380 997.830 ;
        RECT 1066.540 995.700 1071.540 997.830 ;
        RECT 1072.700 995.700 1077.700 997.830 ;
        RECT 1078.860 995.700 1083.860 997.830 ;
        RECT 1085.020 995.700 1090.020 997.830 ;
        RECT 1091.180 995.700 1096.180 997.830 ;
        RECT 1097.340 995.700 1102.340 997.830 ;
        RECT 1103.500 995.700 1108.500 997.830 ;
        RECT 1109.660 995.700 1114.660 997.830 ;
        RECT 1115.820 995.700 1120.820 997.830 ;
        RECT 1121.980 995.700 1126.980 997.830 ;
        RECT 1128.140 995.700 1133.140 997.830 ;
        RECT 1134.300 995.700 1139.300 997.830 ;
        RECT 1140.460 995.700 1145.460 997.830 ;
        RECT 1146.620 995.700 1151.620 997.830 ;
        RECT 1152.780 995.700 1157.780 997.830 ;
        RECT 1158.940 995.700 1163.940 997.830 ;
        RECT 1165.100 995.700 1170.100 997.830 ;
        RECT 1171.260 995.700 1176.260 997.830 ;
        RECT 1177.420 995.700 1182.420 997.830 ;
        RECT 1183.580 995.700 1188.580 997.830 ;
        RECT 1189.740 995.700 1194.740 997.830 ;
        RECT 1195.900 995.700 1200.900 997.830 ;
        RECT 1202.060 995.700 1207.060 997.830 ;
        RECT 1208.220 995.700 1213.220 997.830 ;
        RECT 1214.380 995.700 1219.380 997.830 ;
        RECT 1220.540 995.700 1225.540 997.830 ;
        RECT 1226.700 995.700 1231.700 997.830 ;
        RECT 1232.860 995.700 1237.860 997.830 ;
        RECT 1239.020 995.700 1244.020 997.830 ;
        RECT 1245.180 995.700 1250.180 997.830 ;
        RECT 1251.340 995.700 1256.340 997.830 ;
        RECT 1257.500 995.700 1262.500 997.830 ;
        RECT 1263.660 995.700 1268.660 997.830 ;
        RECT 1269.820 995.700 1274.820 997.830 ;
        RECT 1275.980 995.700 1280.980 997.830 ;
        RECT 1282.140 995.700 1287.140 997.830 ;
        RECT 1288.300 995.700 1293.300 997.830 ;
        RECT 1294.460 995.700 1299.460 997.830 ;
        RECT 1300.620 995.700 1305.620 997.830 ;
        RECT 1306.780 995.700 1311.780 997.830 ;
        RECT 1312.940 995.700 1317.940 997.830 ;
        RECT 1319.100 995.700 1324.100 997.830 ;
        RECT 1325.260 995.700 1330.260 997.830 ;
        RECT 1331.420 995.700 1336.420 997.830 ;
        RECT 1337.580 995.700 1342.580 997.830 ;
        RECT 1343.740 995.700 1348.740 997.830 ;
        RECT 1349.900 995.700 1354.900 997.830 ;
        RECT 1356.060 995.700 1361.060 997.830 ;
        RECT 1362.220 995.700 1367.220 997.830 ;
        RECT 1368.380 995.700 1373.380 997.830 ;
        RECT 1374.540 995.700 1379.540 997.830 ;
        RECT 1380.700 995.700 1385.700 997.830 ;
        RECT 1386.860 995.700 1391.860 997.830 ;
        RECT 1393.020 995.700 1398.020 997.830 ;
        RECT 1399.180 995.700 1404.180 997.830 ;
        RECT 1405.340 995.700 1410.340 997.830 ;
        RECT 1411.500 995.700 1416.500 997.830 ;
        RECT 1417.660 995.700 1422.660 997.830 ;
        RECT 1423.820 995.700 1428.820 997.830 ;
        RECT 1429.980 995.700 1434.980 997.830 ;
        RECT 1436.140 995.700 1441.140 997.830 ;
        RECT 1442.300 995.700 1447.300 997.830 ;
        RECT 1448.460 995.700 1453.460 997.830 ;
        RECT 1454.620 995.700 1459.620 997.830 ;
        RECT 1460.780 995.700 1465.780 997.830 ;
        RECT 1466.940 995.700 1471.940 997.830 ;
        RECT 1473.100 995.700 1478.100 997.830 ;
        RECT 1479.260 995.700 1484.260 997.830 ;
        RECT 1485.420 995.700 1490.420 997.830 ;
        RECT 1491.580 995.700 1496.580 997.830 ;
        RECT 1497.740 995.700 1502.740 997.830 ;
        RECT 1503.900 995.700 1508.900 997.830 ;
        RECT 1510.060 995.700 1515.060 997.830 ;
        RECT 1516.220 995.700 1521.220 997.830 ;
        RECT 1522.380 995.700 1527.380 997.830 ;
        RECT 1528.540 995.700 1533.540 997.830 ;
        RECT 1534.700 995.700 1539.700 997.830 ;
        RECT 1540.860 995.700 1545.860 997.830 ;
        RECT 1547.020 995.700 1552.020 997.830 ;
        RECT 1553.180 995.700 1558.180 997.830 ;
        RECT 1559.340 995.700 1564.340 997.830 ;
        RECT 1565.500 995.700 1570.500 997.830 ;
        RECT 1571.660 995.700 1576.660 997.830 ;
        RECT 1577.820 995.700 1582.820 997.830 ;
        RECT 1583.980 995.700 1588.980 997.830 ;
        RECT 1590.140 995.700 1595.140 997.830 ;
        RECT 1596.300 995.700 1601.300 997.830 ;
        RECT 1602.460 995.700 1607.460 997.830 ;
        RECT 1608.620 995.700 1613.620 997.830 ;
        RECT 1614.780 995.700 1619.780 997.830 ;
        RECT 1620.940 995.700 1625.940 997.830 ;
        RECT 1627.100 995.700 1632.100 997.830 ;
        RECT 1633.260 995.700 1638.260 997.830 ;
        RECT 1639.420 995.700 1644.420 997.830 ;
        RECT 1645.580 995.700 1650.580 997.830 ;
        RECT 1651.740 995.700 1656.740 997.830 ;
        RECT 1657.900 995.700 1662.900 997.830 ;
        RECT 1664.060 995.700 1669.060 997.830 ;
        RECT 1670.220 995.700 1675.220 997.830 ;
        RECT 1676.380 995.700 1681.380 997.830 ;
        RECT 1682.540 995.700 1687.540 997.830 ;
        RECT 1688.700 995.700 1693.700 997.830 ;
        RECT 1694.860 995.700 1699.860 997.830 ;
        RECT 1701.020 995.700 1706.020 997.830 ;
        RECT 1707.180 995.700 1712.180 997.830 ;
        RECT 1713.340 995.700 1718.340 997.830 ;
        RECT 1719.500 995.700 1724.500 997.830 ;
        RECT 1725.660 995.700 1730.660 997.830 ;
        RECT 1731.820 995.700 1790.740 997.830 ;
        RECT 16.380 4.300 1790.740 995.700 ;
        RECT 16.380 0.090 18.740 4.300 ;
        RECT 19.900 0.090 22.100 4.300 ;
        RECT 23.260 0.090 25.460 4.300 ;
        RECT 26.620 0.090 28.820 4.300 ;
        RECT 29.980 0.090 32.180 4.300 ;
        RECT 33.340 0.090 35.540 4.300 ;
        RECT 36.700 0.090 38.900 4.300 ;
        RECT 40.060 0.090 42.260 4.300 ;
        RECT 43.420 0.090 45.620 4.300 ;
        RECT 46.780 0.090 48.980 4.300 ;
        RECT 50.140 0.090 52.340 4.300 ;
        RECT 53.500 0.090 55.700 4.300 ;
        RECT 56.860 0.090 59.060 4.300 ;
        RECT 60.220 0.090 62.420 4.300 ;
        RECT 63.580 0.090 65.780 4.300 ;
        RECT 66.940 0.090 69.140 4.300 ;
        RECT 70.300 0.090 72.500 4.300 ;
        RECT 73.660 0.090 75.860 4.300 ;
        RECT 77.020 0.090 79.220 4.300 ;
        RECT 80.380 0.090 82.580 4.300 ;
        RECT 83.740 0.090 85.940 4.300 ;
        RECT 87.100 0.090 89.300 4.300 ;
        RECT 90.460 0.090 92.660 4.300 ;
        RECT 93.820 0.090 96.020 4.300 ;
        RECT 97.180 0.090 99.380 4.300 ;
        RECT 100.540 0.090 102.740 4.300 ;
        RECT 103.900 0.090 106.100 4.300 ;
        RECT 107.260 0.090 109.460 4.300 ;
        RECT 110.620 0.090 112.820 4.300 ;
        RECT 113.980 0.090 116.180 4.300 ;
        RECT 117.340 0.090 119.540 4.300 ;
        RECT 120.700 0.090 122.900 4.300 ;
        RECT 124.060 0.090 126.260 4.300 ;
        RECT 127.420 0.090 129.620 4.300 ;
        RECT 130.780 0.090 132.980 4.300 ;
        RECT 134.140 0.090 136.340 4.300 ;
        RECT 137.500 0.090 139.700 4.300 ;
        RECT 140.860 0.090 143.060 4.300 ;
        RECT 144.220 0.090 146.420 4.300 ;
        RECT 147.580 0.090 149.780 4.300 ;
        RECT 150.940 0.090 153.140 4.300 ;
        RECT 154.300 0.090 156.500 4.300 ;
        RECT 157.660 0.090 159.860 4.300 ;
        RECT 161.020 0.090 163.220 4.300 ;
        RECT 164.380 0.090 166.580 4.300 ;
        RECT 167.740 0.090 169.940 4.300 ;
        RECT 171.100 0.090 173.300 4.300 ;
        RECT 174.460 0.090 176.660 4.300 ;
        RECT 177.820 0.090 180.020 4.300 ;
        RECT 181.180 0.090 183.380 4.300 ;
        RECT 184.540 0.090 186.740 4.300 ;
        RECT 187.900 0.090 190.100 4.300 ;
        RECT 191.260 0.090 193.460 4.300 ;
        RECT 194.620 0.090 196.820 4.300 ;
        RECT 197.980 0.090 200.180 4.300 ;
        RECT 201.340 0.090 203.540 4.300 ;
        RECT 204.700 0.090 206.900 4.300 ;
        RECT 208.060 0.090 210.260 4.300 ;
        RECT 211.420 0.090 213.620 4.300 ;
        RECT 214.780 0.090 216.980 4.300 ;
        RECT 218.140 0.090 220.340 4.300 ;
        RECT 221.500 0.090 223.700 4.300 ;
        RECT 224.860 0.090 227.060 4.300 ;
        RECT 228.220 0.090 230.420 4.300 ;
        RECT 231.580 0.090 233.780 4.300 ;
        RECT 234.940 0.090 237.140 4.300 ;
        RECT 238.300 0.090 240.500 4.300 ;
        RECT 241.660 0.090 243.860 4.300 ;
        RECT 245.020 0.090 247.220 4.300 ;
        RECT 248.380 0.090 250.580 4.300 ;
        RECT 251.740 0.090 253.940 4.300 ;
        RECT 255.100 0.090 257.300 4.300 ;
        RECT 258.460 0.090 260.660 4.300 ;
        RECT 261.820 0.090 264.020 4.300 ;
        RECT 265.180 0.090 267.380 4.300 ;
        RECT 268.540 0.090 270.740 4.300 ;
        RECT 271.900 0.090 274.100 4.300 ;
        RECT 275.260 0.090 277.460 4.300 ;
        RECT 278.620 0.090 280.820 4.300 ;
        RECT 281.980 0.090 284.180 4.300 ;
        RECT 285.340 0.090 287.540 4.300 ;
        RECT 288.700 0.090 290.900 4.300 ;
        RECT 292.060 0.090 294.260 4.300 ;
        RECT 295.420 0.090 297.620 4.300 ;
        RECT 298.780 0.090 300.980 4.300 ;
        RECT 302.140 0.090 304.340 4.300 ;
        RECT 305.500 0.090 307.700 4.300 ;
        RECT 308.860 0.090 311.060 4.300 ;
        RECT 312.220 0.090 314.420 4.300 ;
        RECT 315.580 0.090 317.780 4.300 ;
        RECT 318.940 0.090 321.140 4.300 ;
        RECT 322.300 0.090 324.500 4.300 ;
        RECT 325.660 0.090 327.860 4.300 ;
        RECT 329.020 0.090 331.220 4.300 ;
        RECT 332.380 0.090 334.580 4.300 ;
        RECT 335.740 0.090 337.940 4.300 ;
        RECT 339.100 0.090 341.300 4.300 ;
        RECT 342.460 0.090 344.660 4.300 ;
        RECT 345.820 0.090 348.020 4.300 ;
        RECT 349.180 0.090 351.380 4.300 ;
        RECT 352.540 0.090 354.740 4.300 ;
        RECT 355.900 0.090 358.100 4.300 ;
        RECT 359.260 0.090 361.460 4.300 ;
        RECT 362.620 0.090 364.820 4.300 ;
        RECT 365.980 0.090 368.180 4.300 ;
        RECT 369.340 0.090 371.540 4.300 ;
        RECT 372.700 0.090 374.900 4.300 ;
        RECT 376.060 0.090 378.260 4.300 ;
        RECT 379.420 0.090 381.620 4.300 ;
        RECT 382.780 0.090 384.980 4.300 ;
        RECT 386.140 0.090 388.340 4.300 ;
        RECT 389.500 0.090 391.700 4.300 ;
        RECT 392.860 0.090 395.060 4.300 ;
        RECT 396.220 0.090 398.420 4.300 ;
        RECT 399.580 0.090 401.780 4.300 ;
        RECT 402.940 0.090 405.140 4.300 ;
        RECT 406.300 0.090 408.500 4.300 ;
        RECT 409.660 0.090 411.860 4.300 ;
        RECT 413.020 0.090 415.220 4.300 ;
        RECT 416.380 0.090 418.580 4.300 ;
        RECT 419.740 0.090 421.940 4.300 ;
        RECT 423.100 0.090 425.300 4.300 ;
        RECT 426.460 0.090 428.660 4.300 ;
        RECT 429.820 0.090 432.020 4.300 ;
        RECT 433.180 0.090 435.380 4.300 ;
        RECT 436.540 0.090 438.740 4.300 ;
        RECT 439.900 0.090 442.100 4.300 ;
        RECT 443.260 0.090 445.460 4.300 ;
        RECT 446.620 0.090 448.820 4.300 ;
        RECT 449.980 0.090 452.180 4.300 ;
        RECT 453.340 0.090 455.540 4.300 ;
        RECT 456.700 0.090 458.900 4.300 ;
        RECT 460.060 0.090 462.260 4.300 ;
        RECT 463.420 0.090 465.620 4.300 ;
        RECT 466.780 0.090 468.980 4.300 ;
        RECT 470.140 0.090 472.340 4.300 ;
        RECT 473.500 0.090 475.700 4.300 ;
        RECT 476.860 0.090 479.060 4.300 ;
        RECT 480.220 0.090 482.420 4.300 ;
        RECT 483.580 0.090 485.780 4.300 ;
        RECT 486.940 0.090 489.140 4.300 ;
        RECT 490.300 0.090 492.500 4.300 ;
        RECT 493.660 0.090 495.860 4.300 ;
        RECT 497.020 0.090 499.220 4.300 ;
        RECT 500.380 0.090 502.580 4.300 ;
        RECT 503.740 0.090 505.940 4.300 ;
        RECT 507.100 0.090 509.300 4.300 ;
        RECT 510.460 0.090 512.660 4.300 ;
        RECT 513.820 0.090 516.020 4.300 ;
        RECT 517.180 0.090 519.380 4.300 ;
        RECT 520.540 0.090 522.740 4.300 ;
        RECT 523.900 0.090 526.100 4.300 ;
        RECT 527.260 0.090 529.460 4.300 ;
        RECT 530.620 0.090 532.820 4.300 ;
        RECT 533.980 0.090 536.180 4.300 ;
        RECT 537.340 0.090 539.540 4.300 ;
        RECT 540.700 0.090 542.900 4.300 ;
        RECT 544.060 0.090 546.260 4.300 ;
        RECT 547.420 0.090 549.620 4.300 ;
        RECT 550.780 0.090 552.980 4.300 ;
        RECT 554.140 0.090 556.340 4.300 ;
        RECT 557.500 0.090 559.700 4.300 ;
        RECT 560.860 0.090 563.060 4.300 ;
        RECT 564.220 0.090 566.420 4.300 ;
        RECT 567.580 0.090 569.780 4.300 ;
        RECT 570.940 0.090 573.140 4.300 ;
        RECT 574.300 0.090 576.500 4.300 ;
        RECT 577.660 0.090 579.860 4.300 ;
        RECT 581.020 0.090 583.220 4.300 ;
        RECT 584.380 0.090 586.580 4.300 ;
        RECT 587.740 0.090 589.940 4.300 ;
        RECT 591.100 0.090 593.300 4.300 ;
        RECT 594.460 0.090 596.660 4.300 ;
        RECT 597.820 0.090 600.020 4.300 ;
        RECT 601.180 0.090 603.380 4.300 ;
        RECT 604.540 0.090 606.740 4.300 ;
        RECT 607.900 0.090 610.100 4.300 ;
        RECT 611.260 0.090 613.460 4.300 ;
        RECT 614.620 0.090 616.820 4.300 ;
        RECT 617.980 0.090 620.180 4.300 ;
        RECT 621.340 0.090 623.540 4.300 ;
        RECT 624.700 0.090 626.900 4.300 ;
        RECT 628.060 0.090 630.260 4.300 ;
        RECT 631.420 0.090 633.620 4.300 ;
        RECT 634.780 0.090 636.980 4.300 ;
        RECT 638.140 0.090 640.340 4.300 ;
        RECT 641.500 0.090 643.700 4.300 ;
        RECT 644.860 0.090 647.060 4.300 ;
        RECT 648.220 0.090 650.420 4.300 ;
        RECT 651.580 0.090 653.780 4.300 ;
        RECT 654.940 0.090 657.140 4.300 ;
        RECT 658.300 0.090 660.500 4.300 ;
        RECT 661.660 0.090 663.860 4.300 ;
        RECT 665.020 0.090 667.220 4.300 ;
        RECT 668.380 0.090 670.580 4.300 ;
        RECT 671.740 0.090 673.940 4.300 ;
        RECT 675.100 0.090 677.300 4.300 ;
        RECT 678.460 0.090 680.660 4.300 ;
        RECT 681.820 0.090 684.020 4.300 ;
        RECT 685.180 0.090 687.380 4.300 ;
        RECT 688.540 0.090 690.740 4.300 ;
        RECT 691.900 0.090 694.100 4.300 ;
        RECT 695.260 0.090 697.460 4.300 ;
        RECT 698.620 0.090 700.820 4.300 ;
        RECT 701.980 0.090 704.180 4.300 ;
        RECT 705.340 0.090 707.540 4.300 ;
        RECT 708.700 0.090 710.900 4.300 ;
        RECT 712.060 0.090 714.260 4.300 ;
        RECT 715.420 0.090 717.620 4.300 ;
        RECT 718.780 0.090 720.980 4.300 ;
        RECT 722.140 0.090 724.340 4.300 ;
        RECT 725.500 0.090 727.700 4.300 ;
        RECT 728.860 0.090 731.060 4.300 ;
        RECT 732.220 0.090 734.420 4.300 ;
        RECT 735.580 0.090 737.780 4.300 ;
        RECT 738.940 0.090 741.140 4.300 ;
        RECT 742.300 0.090 744.500 4.300 ;
        RECT 745.660 0.090 747.860 4.300 ;
        RECT 749.020 0.090 751.220 4.300 ;
        RECT 752.380 0.090 754.580 4.300 ;
        RECT 755.740 0.090 757.940 4.300 ;
        RECT 759.100 0.090 761.300 4.300 ;
        RECT 762.460 0.090 764.660 4.300 ;
        RECT 765.820 0.090 768.020 4.300 ;
        RECT 769.180 0.090 771.380 4.300 ;
        RECT 772.540 0.090 774.740 4.300 ;
        RECT 775.900 0.090 778.100 4.300 ;
        RECT 779.260 0.090 781.460 4.300 ;
        RECT 782.620 0.090 784.820 4.300 ;
        RECT 785.980 0.090 788.180 4.300 ;
        RECT 789.340 0.090 791.540 4.300 ;
        RECT 792.700 0.090 794.900 4.300 ;
        RECT 796.060 0.090 798.260 4.300 ;
        RECT 799.420 0.090 801.620 4.300 ;
        RECT 802.780 0.090 804.980 4.300 ;
        RECT 806.140 0.090 808.340 4.300 ;
        RECT 809.500 0.090 811.700 4.300 ;
        RECT 812.860 0.090 815.060 4.300 ;
        RECT 816.220 0.090 818.420 4.300 ;
        RECT 819.580 0.090 821.780 4.300 ;
        RECT 822.940 0.090 825.140 4.300 ;
        RECT 826.300 0.090 828.500 4.300 ;
        RECT 829.660 0.090 831.860 4.300 ;
        RECT 833.020 0.090 835.220 4.300 ;
        RECT 836.380 0.090 838.580 4.300 ;
        RECT 839.740 0.090 841.940 4.300 ;
        RECT 843.100 0.090 845.300 4.300 ;
        RECT 846.460 0.090 848.660 4.300 ;
        RECT 849.820 0.090 852.020 4.300 ;
        RECT 853.180 0.090 855.380 4.300 ;
        RECT 856.540 0.090 858.740 4.300 ;
        RECT 859.900 0.090 862.100 4.300 ;
        RECT 863.260 0.090 865.460 4.300 ;
        RECT 866.620 0.090 868.820 4.300 ;
        RECT 869.980 0.090 872.180 4.300 ;
        RECT 873.340 0.090 875.540 4.300 ;
        RECT 876.700 0.090 878.900 4.300 ;
        RECT 880.060 0.090 882.260 4.300 ;
        RECT 883.420 0.090 885.620 4.300 ;
        RECT 886.780 0.090 888.980 4.300 ;
        RECT 890.140 0.090 892.340 4.300 ;
        RECT 893.500 0.090 895.700 4.300 ;
        RECT 896.860 0.090 899.060 4.300 ;
        RECT 900.220 0.090 902.420 4.300 ;
        RECT 903.580 0.090 905.780 4.300 ;
        RECT 906.940 0.090 909.140 4.300 ;
        RECT 910.300 0.090 912.500 4.300 ;
        RECT 913.660 0.090 915.860 4.300 ;
        RECT 917.020 0.090 919.220 4.300 ;
        RECT 920.380 0.090 922.580 4.300 ;
        RECT 923.740 0.090 925.940 4.300 ;
        RECT 927.100 0.090 929.300 4.300 ;
        RECT 930.460 0.090 932.660 4.300 ;
        RECT 933.820 0.090 936.020 4.300 ;
        RECT 937.180 0.090 939.380 4.300 ;
        RECT 940.540 0.090 942.740 4.300 ;
        RECT 943.900 0.090 946.100 4.300 ;
        RECT 947.260 0.090 949.460 4.300 ;
        RECT 950.620 0.090 952.820 4.300 ;
        RECT 953.980 0.090 956.180 4.300 ;
        RECT 957.340 0.090 959.540 4.300 ;
        RECT 960.700 0.090 962.900 4.300 ;
        RECT 964.060 0.090 966.260 4.300 ;
        RECT 967.420 0.090 969.620 4.300 ;
        RECT 970.780 0.090 972.980 4.300 ;
        RECT 974.140 0.090 976.340 4.300 ;
        RECT 977.500 0.090 979.700 4.300 ;
        RECT 980.860 0.090 983.060 4.300 ;
        RECT 984.220 0.090 986.420 4.300 ;
        RECT 987.580 0.090 989.780 4.300 ;
        RECT 990.940 0.090 993.140 4.300 ;
        RECT 994.300 0.090 996.500 4.300 ;
        RECT 997.660 0.090 999.860 4.300 ;
        RECT 1001.020 0.090 1003.220 4.300 ;
        RECT 1004.380 0.090 1006.580 4.300 ;
        RECT 1007.740 0.090 1009.940 4.300 ;
        RECT 1011.100 0.090 1013.300 4.300 ;
        RECT 1014.460 0.090 1016.660 4.300 ;
        RECT 1017.820 0.090 1020.020 4.300 ;
        RECT 1021.180 0.090 1023.380 4.300 ;
        RECT 1024.540 0.090 1026.740 4.300 ;
        RECT 1027.900 0.090 1030.100 4.300 ;
        RECT 1031.260 0.090 1033.460 4.300 ;
        RECT 1034.620 0.090 1036.820 4.300 ;
        RECT 1037.980 0.090 1040.180 4.300 ;
        RECT 1041.340 0.090 1043.540 4.300 ;
        RECT 1044.700 0.090 1046.900 4.300 ;
        RECT 1048.060 0.090 1050.260 4.300 ;
        RECT 1051.420 0.090 1053.620 4.300 ;
        RECT 1054.780 0.090 1056.980 4.300 ;
        RECT 1058.140 0.090 1060.340 4.300 ;
        RECT 1061.500 0.090 1063.700 4.300 ;
        RECT 1064.860 0.090 1067.060 4.300 ;
        RECT 1068.220 0.090 1070.420 4.300 ;
        RECT 1071.580 0.090 1073.780 4.300 ;
        RECT 1074.940 0.090 1077.140 4.300 ;
        RECT 1078.300 0.090 1080.500 4.300 ;
        RECT 1081.660 0.090 1083.860 4.300 ;
        RECT 1085.020 0.090 1087.220 4.300 ;
        RECT 1088.380 0.090 1090.580 4.300 ;
        RECT 1091.740 0.090 1093.940 4.300 ;
        RECT 1095.100 0.090 1097.300 4.300 ;
        RECT 1098.460 0.090 1100.660 4.300 ;
        RECT 1101.820 0.090 1104.020 4.300 ;
        RECT 1105.180 0.090 1107.380 4.300 ;
        RECT 1108.540 0.090 1110.740 4.300 ;
        RECT 1111.900 0.090 1114.100 4.300 ;
        RECT 1115.260 0.090 1117.460 4.300 ;
        RECT 1118.620 0.090 1120.820 4.300 ;
        RECT 1121.980 0.090 1124.180 4.300 ;
        RECT 1125.340 0.090 1127.540 4.300 ;
        RECT 1128.700 0.090 1130.900 4.300 ;
        RECT 1132.060 0.090 1134.260 4.300 ;
        RECT 1135.420 0.090 1137.620 4.300 ;
        RECT 1138.780 0.090 1140.980 4.300 ;
        RECT 1142.140 0.090 1144.340 4.300 ;
        RECT 1145.500 0.090 1147.700 4.300 ;
        RECT 1148.860 0.090 1151.060 4.300 ;
        RECT 1152.220 0.090 1154.420 4.300 ;
        RECT 1155.580 0.090 1157.780 4.300 ;
        RECT 1158.940 0.090 1161.140 4.300 ;
        RECT 1162.300 0.090 1164.500 4.300 ;
        RECT 1165.660 0.090 1167.860 4.300 ;
        RECT 1169.020 0.090 1171.220 4.300 ;
        RECT 1172.380 0.090 1174.580 4.300 ;
        RECT 1175.740 0.090 1177.940 4.300 ;
        RECT 1179.100 0.090 1181.300 4.300 ;
        RECT 1182.460 0.090 1184.660 4.300 ;
        RECT 1185.820 0.090 1188.020 4.300 ;
        RECT 1189.180 0.090 1191.380 4.300 ;
        RECT 1192.540 0.090 1194.740 4.300 ;
        RECT 1195.900 0.090 1198.100 4.300 ;
        RECT 1199.260 0.090 1201.460 4.300 ;
        RECT 1202.620 0.090 1204.820 4.300 ;
        RECT 1205.980 0.090 1208.180 4.300 ;
        RECT 1209.340 0.090 1211.540 4.300 ;
        RECT 1212.700 0.090 1214.900 4.300 ;
        RECT 1216.060 0.090 1218.260 4.300 ;
        RECT 1219.420 0.090 1221.620 4.300 ;
        RECT 1222.780 0.090 1224.980 4.300 ;
        RECT 1226.140 0.090 1228.340 4.300 ;
        RECT 1229.500 0.090 1231.700 4.300 ;
        RECT 1232.860 0.090 1235.060 4.300 ;
        RECT 1236.220 0.090 1238.420 4.300 ;
        RECT 1239.580 0.090 1241.780 4.300 ;
        RECT 1242.940 0.090 1245.140 4.300 ;
        RECT 1246.300 0.090 1248.500 4.300 ;
        RECT 1249.660 0.090 1251.860 4.300 ;
        RECT 1253.020 0.090 1255.220 4.300 ;
        RECT 1256.380 0.090 1258.580 4.300 ;
        RECT 1259.740 0.090 1261.940 4.300 ;
        RECT 1263.100 0.090 1265.300 4.300 ;
        RECT 1266.460 0.090 1268.660 4.300 ;
        RECT 1269.820 0.090 1272.020 4.300 ;
        RECT 1273.180 0.090 1275.380 4.300 ;
        RECT 1276.540 0.090 1278.740 4.300 ;
        RECT 1279.900 0.090 1282.100 4.300 ;
        RECT 1283.260 0.090 1285.460 4.300 ;
        RECT 1286.620 0.090 1288.820 4.300 ;
        RECT 1289.980 0.090 1292.180 4.300 ;
        RECT 1293.340 0.090 1295.540 4.300 ;
        RECT 1296.700 0.090 1298.900 4.300 ;
        RECT 1300.060 0.090 1302.260 4.300 ;
        RECT 1303.420 0.090 1305.620 4.300 ;
        RECT 1306.780 0.090 1308.980 4.300 ;
        RECT 1310.140 0.090 1312.340 4.300 ;
        RECT 1313.500 0.090 1315.700 4.300 ;
        RECT 1316.860 0.090 1319.060 4.300 ;
        RECT 1320.220 0.090 1322.420 4.300 ;
        RECT 1323.580 0.090 1325.780 4.300 ;
        RECT 1326.940 0.090 1329.140 4.300 ;
        RECT 1330.300 0.090 1332.500 4.300 ;
        RECT 1333.660 0.090 1335.860 4.300 ;
        RECT 1337.020 0.090 1339.220 4.300 ;
        RECT 1340.380 0.090 1342.580 4.300 ;
        RECT 1343.740 0.090 1345.940 4.300 ;
        RECT 1347.100 0.090 1349.300 4.300 ;
        RECT 1350.460 0.090 1352.660 4.300 ;
        RECT 1353.820 0.090 1356.020 4.300 ;
        RECT 1357.180 0.090 1359.380 4.300 ;
        RECT 1360.540 0.090 1362.740 4.300 ;
        RECT 1363.900 0.090 1366.100 4.300 ;
        RECT 1367.260 0.090 1369.460 4.300 ;
        RECT 1370.620 0.090 1372.820 4.300 ;
        RECT 1373.980 0.090 1376.180 4.300 ;
        RECT 1377.340 0.090 1379.540 4.300 ;
        RECT 1380.700 0.090 1382.900 4.300 ;
        RECT 1384.060 0.090 1386.260 4.300 ;
        RECT 1387.420 0.090 1389.620 4.300 ;
        RECT 1390.780 0.090 1392.980 4.300 ;
        RECT 1394.140 0.090 1396.340 4.300 ;
        RECT 1397.500 0.090 1399.700 4.300 ;
        RECT 1400.860 0.090 1403.060 4.300 ;
        RECT 1404.220 0.090 1406.420 4.300 ;
        RECT 1407.580 0.090 1409.780 4.300 ;
        RECT 1410.940 0.090 1413.140 4.300 ;
        RECT 1414.300 0.090 1416.500 4.300 ;
        RECT 1417.660 0.090 1419.860 4.300 ;
        RECT 1421.020 0.090 1423.220 4.300 ;
        RECT 1424.380 0.090 1426.580 4.300 ;
        RECT 1427.740 0.090 1429.940 4.300 ;
        RECT 1431.100 0.090 1433.300 4.300 ;
        RECT 1434.460 0.090 1436.660 4.300 ;
        RECT 1437.820 0.090 1440.020 4.300 ;
        RECT 1441.180 0.090 1443.380 4.300 ;
        RECT 1444.540 0.090 1446.740 4.300 ;
        RECT 1447.900 0.090 1450.100 4.300 ;
        RECT 1451.260 0.090 1453.460 4.300 ;
        RECT 1454.620 0.090 1456.820 4.300 ;
        RECT 1457.980 0.090 1460.180 4.300 ;
        RECT 1461.340 0.090 1463.540 4.300 ;
        RECT 1464.700 0.090 1466.900 4.300 ;
        RECT 1468.060 0.090 1470.260 4.300 ;
        RECT 1471.420 0.090 1473.620 4.300 ;
        RECT 1474.780 0.090 1476.980 4.300 ;
        RECT 1478.140 0.090 1480.340 4.300 ;
        RECT 1481.500 0.090 1483.700 4.300 ;
        RECT 1484.860 0.090 1487.060 4.300 ;
        RECT 1488.220 0.090 1490.420 4.300 ;
        RECT 1491.580 0.090 1493.780 4.300 ;
        RECT 1494.940 0.090 1497.140 4.300 ;
        RECT 1498.300 0.090 1500.500 4.300 ;
        RECT 1501.660 0.090 1503.860 4.300 ;
        RECT 1505.020 0.090 1507.220 4.300 ;
        RECT 1508.380 0.090 1510.580 4.300 ;
        RECT 1511.740 0.090 1513.940 4.300 ;
        RECT 1515.100 0.090 1517.300 4.300 ;
        RECT 1518.460 0.090 1520.660 4.300 ;
        RECT 1521.820 0.090 1524.020 4.300 ;
        RECT 1525.180 0.090 1527.380 4.300 ;
        RECT 1528.540 0.090 1530.740 4.300 ;
        RECT 1531.900 0.090 1534.100 4.300 ;
        RECT 1535.260 0.090 1537.460 4.300 ;
        RECT 1538.620 0.090 1540.820 4.300 ;
        RECT 1541.980 0.090 1544.180 4.300 ;
        RECT 1545.340 0.090 1547.540 4.300 ;
        RECT 1548.700 0.090 1550.900 4.300 ;
        RECT 1552.060 0.090 1554.260 4.300 ;
        RECT 1555.420 0.090 1557.620 4.300 ;
        RECT 1558.780 0.090 1560.980 4.300 ;
        RECT 1562.140 0.090 1564.340 4.300 ;
        RECT 1565.500 0.090 1567.700 4.300 ;
        RECT 1568.860 0.090 1571.060 4.300 ;
        RECT 1572.220 0.090 1574.420 4.300 ;
        RECT 1575.580 0.090 1577.780 4.300 ;
        RECT 1578.940 0.090 1581.140 4.300 ;
        RECT 1582.300 0.090 1584.500 4.300 ;
        RECT 1585.660 0.090 1587.860 4.300 ;
        RECT 1589.020 0.090 1591.220 4.300 ;
        RECT 1592.380 0.090 1594.580 4.300 ;
        RECT 1595.740 0.090 1597.940 4.300 ;
        RECT 1599.100 0.090 1601.300 4.300 ;
        RECT 1602.460 0.090 1604.660 4.300 ;
        RECT 1605.820 0.090 1608.020 4.300 ;
        RECT 1609.180 0.090 1611.380 4.300 ;
        RECT 1612.540 0.090 1614.740 4.300 ;
        RECT 1615.900 0.090 1618.100 4.300 ;
        RECT 1619.260 0.090 1621.460 4.300 ;
        RECT 1622.620 0.090 1624.820 4.300 ;
        RECT 1625.980 0.090 1628.180 4.300 ;
        RECT 1629.340 0.090 1631.540 4.300 ;
        RECT 1632.700 0.090 1634.900 4.300 ;
        RECT 1636.060 0.090 1638.260 4.300 ;
        RECT 1639.420 0.090 1641.620 4.300 ;
        RECT 1642.780 0.090 1644.980 4.300 ;
        RECT 1646.140 0.090 1648.340 4.300 ;
        RECT 1649.500 0.090 1651.700 4.300 ;
        RECT 1652.860 0.090 1655.060 4.300 ;
        RECT 1656.220 0.090 1658.420 4.300 ;
        RECT 1659.580 0.090 1661.780 4.300 ;
        RECT 1662.940 0.090 1665.140 4.300 ;
        RECT 1666.300 0.090 1668.500 4.300 ;
        RECT 1669.660 0.090 1671.860 4.300 ;
        RECT 1673.020 0.090 1675.220 4.300 ;
        RECT 1676.380 0.090 1678.580 4.300 ;
        RECT 1679.740 0.090 1681.940 4.300 ;
        RECT 1683.100 0.090 1685.300 4.300 ;
        RECT 1686.460 0.090 1688.660 4.300 ;
        RECT 1689.820 0.090 1692.020 4.300 ;
        RECT 1693.180 0.090 1695.380 4.300 ;
        RECT 1696.540 0.090 1698.740 4.300 ;
        RECT 1699.900 0.090 1702.100 4.300 ;
        RECT 1703.260 0.090 1705.460 4.300 ;
        RECT 1706.620 0.090 1708.820 4.300 ;
        RECT 1709.980 0.090 1712.180 4.300 ;
        RECT 1713.340 0.090 1715.540 4.300 ;
        RECT 1716.700 0.090 1718.900 4.300 ;
        RECT 1720.060 0.090 1722.260 4.300 ;
        RECT 1723.420 0.090 1725.620 4.300 ;
        RECT 1726.780 0.090 1728.980 4.300 ;
        RECT 1730.140 0.090 1732.340 4.300 ;
        RECT 1733.500 0.090 1735.700 4.300 ;
        RECT 1736.860 0.090 1739.060 4.300 ;
        RECT 1740.220 0.090 1742.420 4.300 ;
        RECT 1743.580 0.090 1745.780 4.300 ;
        RECT 1746.940 0.090 1749.140 4.300 ;
        RECT 1750.300 0.090 1752.500 4.300 ;
        RECT 1753.660 0.090 1755.860 4.300 ;
        RECT 1757.020 0.090 1759.220 4.300 ;
        RECT 1760.380 0.090 1762.580 4.300 ;
        RECT 1763.740 0.090 1765.940 4.300 ;
        RECT 1767.100 0.090 1769.300 4.300 ;
        RECT 1770.460 0.090 1772.660 4.300 ;
        RECT 1773.820 0.090 1776.020 4.300 ;
        RECT 1777.180 0.090 1779.380 4.300 ;
        RECT 1780.540 0.090 1790.740 4.300 ;
      LAYER Metal3 ;
        RECT 16.330 0.140 1790.790 997.780 ;
      LAYER Metal4 ;
        RECT 159.740 984.520 1376.900 994.470 ;
        RECT 159.740 26.410 175.540 984.520 ;
        RECT 177.740 26.410 252.340 984.520 ;
        RECT 254.540 26.410 329.140 984.520 ;
        RECT 331.340 26.410 405.940 984.520 ;
        RECT 408.140 26.410 482.740 984.520 ;
        RECT 484.940 26.410 559.540 984.520 ;
        RECT 561.740 26.410 636.340 984.520 ;
        RECT 638.540 26.410 713.140 984.520 ;
        RECT 715.340 26.410 789.940 984.520 ;
        RECT 792.140 26.410 866.740 984.520 ;
        RECT 868.940 26.410 943.540 984.520 ;
        RECT 945.740 26.410 1020.340 984.520 ;
        RECT 1022.540 26.410 1097.140 984.520 ;
        RECT 1099.340 26.410 1173.940 984.520 ;
        RECT 1176.140 26.410 1250.740 984.520 ;
        RECT 1252.940 26.410 1327.540 984.520 ;
        RECT 1329.740 26.410 1376.900 984.520 ;
  END
END io_interface
END LIBRARY

