* NGSPICE file created from io_interface.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

.subckt io_interface Serial_input Serial_output analog_io[0] analog_io[10] analog_io[11]
+ analog_io[12] analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17]
+ analog_io[18] analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22]
+ analog_io[23] analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28]
+ analog_io[2] analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8]
+ analog_io[9] clk data_mem_addr[0] data_mem_addr[1] data_mem_addr[2] data_mem_addr[3]
+ data_mem_addr[4] data_mem_addr[5] data_mem_addr[6] data_mem_addr[7] data_mem_sel
+ data_read_data[0] data_read_data[10] data_read_data[11] data_read_data[12] data_read_data[13]
+ data_read_data[14] data_read_data[15] data_read_data[1] data_read_data[2] data_read_data[3]
+ data_read_data[4] data_read_data[5] data_read_data[6] data_read_data[7] data_read_data[8]
+ data_read_data[9] data_write_data[0] data_write_data[10] data_write_data[11] data_write_data[12]
+ data_write_data[13] data_write_data[14] data_write_data[15] data_write_data[1] data_write_data[2]
+ data_write_data[3] data_write_data[4] data_write_data[5] data_write_data[6] data_write_data[7]
+ data_write_data[8] data_write_data[9] dataw_en dataw_en_8bit[0] dataw_en_8bit[1]
+ dataw_en_8bit[2] dataw_en_8bit[3] dataw_en_8bit[4] dataw_en_8bit[5] dataw_en_8bit[6]
+ dataw_en_8bit[7] hlt instr[0] instr[10] instr[11] instr[12] instr[13] instr[14]
+ instr[15] instr[1] instr[2] instr[3] instr[4] instr[5] instr[6] instr[7] instr[8]
+ instr[9] instr_mem_addr[0] instr_mem_addr[1] instr_mem_addr[2] instr_mem_addr[3]
+ instr_mem_addr[4] instr_mem_addr[5] instr_mem_addr[6] instr_mem_addr[7] instr_mem_sel
+ instr_write_data[0] instr_write_data[10] instr_write_data[11] instr_write_data[12]
+ instr_write_data[13] instr_write_data[14] instr_write_data[15] instr_write_data[1]
+ instr_write_data[2] instr_write_data[3] instr_write_data[4] instr_write_data[5]
+ instr_write_data[6] instr_write_data[7] instr_write_data[8] instr_write_data[9]
+ instrw_en instrw_en_8bit[0] instrw_en_8bit[1] instrw_en_8bit[2] instrw_en_8bit[3]
+ instrw_en_8bit[4] instrw_en_8bit[5] instrw_en_8bit[6] instrw_en_8bit[7] io_in[0]
+ io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] irq[0] irq[1] irq[2]
+ la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101]
+ la_oenb[102] la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108]
+ la_oenb[109] la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114]
+ la_oenb[115] la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120]
+ la_oenb[121] la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18]
+ la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24]
+ la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30]
+ la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4]
+ la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62]
+ la_oenb[63] la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69]
+ la_oenb[6] la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75]
+ la_oenb[76] la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81]
+ la_oenb[82] la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88]
+ la_oenb[89] la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94]
+ la_oenb[95] la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] reset start
+ uP_data_mem_addr[0] uP_data_mem_addr[1] uP_data_mem_addr[2] uP_data_mem_addr[3]
+ uP_data_mem_addr[4] uP_data_mem_addr[5] uP_data_mem_addr[6] uP_data_mem_addr[7]
+ uP_dataw_en uP_instr[0] uP_instr[10] uP_instr[11] uP_instr[12] uP_instr[13] uP_instr[14]
+ uP_instr[15] uP_instr[1] uP_instr[2] uP_instr[3] uP_instr[4] uP_instr[5] uP_instr[6]
+ uP_instr[7] uP_instr[8] uP_instr[9] uP_instr_mem_addr[0] uP_instr_mem_addr[10] uP_instr_mem_addr[11]
+ uP_instr_mem_addr[12] uP_instr_mem_addr[1] uP_instr_mem_addr[2] uP_instr_mem_addr[3]
+ uP_instr_mem_addr[4] uP_instr_mem_addr[5] uP_instr_mem_addr[6] uP_instr_mem_addr[7]
+ uP_instr_mem_addr[8] uP_instr_mem_addr[9] uP_write_data[0] uP_write_data[10] uP_write_data[11]
+ uP_write_data[12] uP_write_data[13] uP_write_data[14] uP_write_data[15] uP_write_data[1]
+ uP_write_data[2] uP_write_data[3] uP_write_data[4] uP_write_data[5] uP_write_data[6]
+ uP_write_data[7] uP_write_data[8] uP_write_data[9] vdd vss wb_clk_i wb_rst_i wbs_ack_o
+ wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_116_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input108_I la_data_in[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input73_I la_data_in[117] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_8917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0496__A2 net699 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_196_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0559__I0 _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_220_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0985_ _0164_ _0096_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput423 net423 data_mem_addr[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput434 net434 data_write_data[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput445 net445 dataw_en_8bit[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput456 net456 instr_mem_addr[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_64_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput467 net467 instr_write_data[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput478 net478 instrw_en_8bit[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput489 net489 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_5_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input225_I la_oenb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0961__I0 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout683 net684 net683 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_150_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout694 net53 net694 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_76_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_210_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0770_ _0393_ net555 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_239_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0952__I0 net695 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1253_ net396 net663 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_204_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1184_ net358 analog_io[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_209_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0968_ _0086_ net523 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0899_ _0047_ net617 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_7309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input175_I la_data_in[94] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input342_I wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input36_I io_in[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0943__I0 net699 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_9212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_8577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_8599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0836__I _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0822_ _0422_ net581 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0753_ net632 net105 _0382_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0473__S1 _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0684_ _0321_ _0342_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1236_ net378 net645 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1167_ net371 analog_io[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0605__A2 net694 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0481__I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input292_I la_oenb[85] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1030__A2 _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_240_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_238_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_7695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1021_ _0124_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0805_ net438 net130 _0409_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1012__A2 _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0736_ net640 net97 _0371_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0667_ _0322_ _0323_ _0324_ _0325_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_135_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0598_ _0277_ net630 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input138_I la_data_in[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0476__I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1219_ net687 net478 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input305_I la_oenb[97] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput301 la_oenb[93] net301 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput312 uP_data_mem_addr[3] net312 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_6268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput323 uP_instr_mem_addr[5] net323 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_6279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput334 uP_write_data[2] net334 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_195_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0514__A1 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput345 wbs_adr_i[10] net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_721 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__0514__B2 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput356 wbs_adr_i[20] net356 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_732 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput367 wbs_adr_i[30] net367 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_743 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_236_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput378 wbs_dat_i[10] net378 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput389 wbs_dat_i[20] net389 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xio_interface_754 irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_91_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_765 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_166_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_776 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_75_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_224_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1010__I _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0521_ _0201_ net49 _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_177_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0452_ _0173_ _0174_ _0171_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_234_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0505__A1 instr_load_addr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0505__B2 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1004_ _0187_ _0107_ instr_load_addr\[5\] _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_147_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0992__A1 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0719_ _0364_ net532 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_10971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input255_I la_oenb[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_218_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_208_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_output641_I net641 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput120 la_data_in[44] net120 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput131 la_data_in[54] net131 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput142 la_data_in[64] net142 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput153 la_data_in[74] net153 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput164 la_data_in[84] net164 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_20_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput175 la_data_in[94] net175 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_79_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput186 la_oenb[104] net186 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput197 la_oenb[114] net197 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_103_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_10223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput605 net605 la_data_out[82] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput616 net616 la_data_out[92] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput627 net627 uP_instr[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput638 net638 uP_instr[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput649 net649 wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_29_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0504_ _0201_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_136_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_231_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_241_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input372_I wbs_adr_i[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input66_I la_data_in[110] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_11480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_199_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0984_ _0094_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_207_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput424 net424 data_write_data[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_233_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput435 net435 data_write_data[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput446 net446 dataw_en_8bit[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput457 net457 instr_write_data[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput468 net468 instr_write_data[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput479 net479 instrw_en_8bit[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_236_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input120_I la_data_in[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input218_I la_oenb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_8759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_215_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output437_I net437 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0961__I1 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout684 net685 net684 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout695 net46 net695 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_41_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1252_ net395 net662 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_238_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1183_ net357 analog_io[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0468__I0 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_200_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0967_ net693 net79 _0085_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0898_ net497 net174 _0043_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__0640__I0 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input168_I la_data_in[88] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input335_I uP_write_data[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input29_I instr[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0459__I0 _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0821_ net430 net138 _0419_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0752_ _0383_ net546 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0683_ _0326_ _0331_ _0336_ _0341_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_100_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_215_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1235_ net408 net675 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1166_ net370 analog_io[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_4_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0861__I0 net416 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input285_I la_oenb[79] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0937__I _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_229_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_240_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_240_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0852__I0 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_200_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_9076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1020_ _0123_ net699 _0109_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0843__I0 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0804_ _0412_ net572 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0735_ _0373_ net539 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_219_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0666_ net230 net229 net233 net232 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_67_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0597_ net21 _0273_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_230_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_217_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1218_ net688 net477 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0693__S _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input200_I la_oenb[117] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input96_I la_data_in[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0834__I0 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput302 la_oenb[94] net302 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput313 uP_data_mem_addr[4] net313 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_6269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput324 uP_instr_mem_addr[6] net324 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_233_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput335 uP_write_data[3] net335 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_209_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0514__A2 _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput346 wbs_adr_i[11] net346 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_5557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_722 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_5_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput357 wbs_adr_i[21] net357 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_733 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput368 wbs_adr_i[31] net368 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_744 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_188_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput379 wbs_dat_i[11] net379 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_755 irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_766 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_2_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_777 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_131_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0520_ net7 _0223_ _0224_ net24 _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_171_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0451_ net8 net25 data_load_addr\[1\] instr_load_addr\[1\] _0166_ _0168_ _0174_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_7460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1003_ _0110_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1201__I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_206_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0718_ net88 _0345_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_63_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0649_ net279 net278 net281 net280 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_24_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input150_I la_data_in[71] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input248_I la_oenb[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_210_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input11_I data_read_data[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output467_I net467 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output634_I net634 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_6044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput110 la_data_in[35] net110 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_6077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput121 la_data_in[45] net121 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput132 la_data_in[55] net132 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput143 la_data_in[65] net143 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_79_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput154 la_data_in[75] net154 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput165 la_data_in[85] net165 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_59_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput176 la_data_in[95] net176 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput187 la_oenb[105] net187 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput198 la_oenb[115] net198 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_105_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput606 net606 la_data_out[83] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput617 net617 la_data_out[93] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput628 net628 uP_instr[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_236_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput639 net639 uP_instr[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0503_ _0202_ _0215_ _0216_ net483 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_193_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input3_I data_read_data[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0971__S _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_225_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input198_I la_oenb[115] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input365_I wbs_adr_i[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input59_I la_data_in[104] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1016__I _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0983_ _0094_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0590__I _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_218_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput425 net425 data_write_data[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput436 net436 data_write_data[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput447 net447 dataw_en_8bit[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput458 net458 instr_write_data[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput469 net469 instr_write_data[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input113_I la_data_in[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_244_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1060__A1 _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout685 net686 net685 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_219_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout696 net45 net696 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1051__A1 data_load_addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_196_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0786__S _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1251_ net394 net661 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_215_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_209_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1182_ net356 analog_io[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_228_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0468__I1 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0966_ _0069_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_119_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1042__A1 _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0897_ _0046_ net616 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input230_I la_oenb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input328_I uP_write_data[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0495__I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1033__A1 _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_245_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0820_ _0421_ net579 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1024__A1 _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0458__S0 _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0751_ net631 net103 _0382_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0682_ _0337_ _0338_ _0339_ _0340_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_9770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1234_ net407 net674 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1165_ net369 analog_io[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_20_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1204__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0949_ _0076_ net514 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input180_I la_data_in[99] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input278_I la_oenb[72] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input41_I io_in[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output497_I net497 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1006__A1 _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0517__B1 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0540__I0 _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0863__I _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0803_ net437 net129 _0409_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0734_ net639 net96 _0371_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout695_I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0665_ net226 net225 net228 net227 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_154_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0596_ _0276_ net629 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1020__I1 net699 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1217_ net689 net476 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1079_ _0016_ net702 net678 instr_load_addr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_181_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input395_I wbs_dat_i[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input89_I la_data_in[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput303 la_oenb[95] net303 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput314 uP_data_mem_addr[5] net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput325 uP_instr_mem_addr[7] net325 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput336 uP_write_data[4] net336 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_712 Serial_output vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput347 wbs_adr_i[12] net347 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_723 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput358 wbs_adr_i[22] net358 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_734 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_233_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput369 wbs_adr_i[3] net369 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xio_interface_745 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_229_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_756 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_79_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_767 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_4868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_778 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_4879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_207_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0450_ net35 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_216_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1002__I1 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0794__S _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1002_ _0108_ _0186_ _0109_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_169_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout708_I net709 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0969__S _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0717_ _0363_ net531 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0648_ net270 net269 net272 net271 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_28_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0768__I _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0579_ net28 _0260_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_230_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input143_I la_data_in[65] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input310_I uP_data_mem_addr[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input408_I wbs_dat_i[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_213_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output627_I net627 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput100 la_data_in[26] net100 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput111 la_data_in[36] net111 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput122 la_data_in[46] net122 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput133 la_data_in[56] net133 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0499__A2 net698 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput144 la_data_in[66] net144 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_24_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput155 la_data_in[76] net155 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput166 la_data_in[86] net166 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput177 la_data_in[96] net177 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_40_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput188 la_oenb[106] net188 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_3920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput199 la_oenb[116] net199 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_2_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_220_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_103_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput607 net607 la_data_out[84] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput618 net618 la_data_out[94] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput629 net629 uP_instr[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_218_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0502_ _0211_ net697 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_7291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0734__I0 net639 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1212__I net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0662__A2 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input260_I la_oenb[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input358_I wbs_adr_i[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0973__I0 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0725__I0 net635 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0982_ _0093_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput415 net686 clk vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput426 net426 data_write_data[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput437 net437 data_write_data[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput448 net448 dataw_en_8bit[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_10077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput459 net459 instr_write_data[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1207__I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input106_I la_data_in[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input71_I la_data_in[115] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_8717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0571__A1 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout686 net415 net686 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_150_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0956__I _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout697 net44 net697 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1250_ net393 net660 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1181_ net354 analog_io[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0468__I2 data_load_addr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0965_ _0084_ net522 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1042__A2 _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0896_ net496 net173 _0043_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0977__S _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input223_I la_oenb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0686__I _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_235_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0750_ _0376_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__0458__S1 _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0681_ net248 net247 net250 net249 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_48_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_234_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1233_ net406 net673 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1164_ net366 analog_io[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_98_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1015__A2 instr_load_addr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0948_ net697 net70 _0075_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_198_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0879_ _0036_ net607 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input173_I la_data_in[92] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input340_I uP_write_data[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input34_I io_in[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_9012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0517__A1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0517__B2 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_212_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0540__I1 net314 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1040__I _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0802_ _0411_ net571 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0733_ _0372_ net538 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0664_ net217 net216 net219 net218 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_171_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0595_ net20 _0273_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1215__I net690 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1216_ net690 net475 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1078_ _0015_ net705 net678 instr_load_addr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_146_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0995__A1 instr_load_addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input290_I la_oenb[83] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input388_I wbs_dat_i[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_235_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput304 la_oenb[96] net304 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput315 uP_data_mem_addr[6] net315 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_216_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput326 uP_write_data[0] net326 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput337 uP_write_data[5] net337 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_713 data_mem_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_152_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput348 wbs_adr_i[13] net348 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_724 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_5_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput359 wbs_adr_i[23] net359 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_735 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_746 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_757 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xio_interface_768 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_4869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_243_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_107_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0986__A1 _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1001_ _0093_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_212_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0716_ net87 _0345_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0647_ net274 net273 net277 net276 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_236_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0578_ _0266_ net636 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_217_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input136_I la_data_in[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input303_I la_oenb[95] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput101 la_data_in[27] net101 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_172_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput112 la_data_in[37] net112 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output522_I net522 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput123 la_data_in[47] net123 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput134 la_data_in[57] net134 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput145 la_data_in[67] net145 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput156 la_data_in[77] net156 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_131_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput167 la_data_in[87] net167 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput178 la_data_in[97] net178 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_44_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput189 la_oenb[107] net189 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_3910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_103_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_207_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput608 net608 la_data_out[85] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput619 net619 la_data_out[95] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_233_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0501_ instr_load_addr\[10\] _0204_ _0206_ net2 _0209_ net19 _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_138_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0662__A3 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input253_I la_oenb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_159_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0964__I1 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0981_ _0203_ _0281_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_35_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput416 net416 data_mem_addr[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput427 net427 data_write_data[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__0599__I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput438 net438 data_write_data[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_173_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput449 net449 instr_mem_addr[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1223__I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_224_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input370_I wbs_adr_i[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_8707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input64_I la_data_in[109] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_11280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout676 net677 net676 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout687 net688 net687 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_189_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout698 net43 net698 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_41_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_230_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0634__I0 net695 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1180_ net353 analog_io[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_65_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_220_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0882__I _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0468__I3 _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0964_ net687 net78 _0080_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_242_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0625__I0 net699 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0895_ _0045_ net615 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input216_I la_oenb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0616__I0 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output435_I net435 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0855__I0 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0607__I0 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0680_ net244 net243 net246 net245 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_139_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1232_ net405 net672 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1163_ net355 analog_io[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_96_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1094_ _0007_ net707 net682 data_load_addr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_228_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0846__I0 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1015__A3 _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0947_ _0069_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0878_ net423 net164 _0033_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input166_I la_data_in[86] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input333_I uP_write_data[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input27_I instr[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0837__I0 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0517__A2 _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0697__I _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0828__I0 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0801_ net436 net128 _0409_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0732_ net638 net95 _0371_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0663_ net222 net221 net224 net223 _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_9580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0594_ _0275_ net628 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_174_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_187_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1215_ net690 net474 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1077_ _0014_ net700 net677 instr_load_addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_213_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0819__I0 net429 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0995__A2 _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input283_I la_oenb[77] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput305 la_oenb[97] net305 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_40_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput316 uP_data_mem_addr[7] net316 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput327 uP_write_data[10] net327 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_44_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput338 uP_write_data[6] net338 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_118_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_714 instr_mem_sel vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput349 wbs_adr_i[14] net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_725 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_736 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_2_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_747 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_217_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_758 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_211_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_769 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_166_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0683__A1 _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_224_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_223_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0986__A2 _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1000_ _0187_ _0107_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0715_ _0362_ net530 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_10942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0646_ _0301_ _0302_ _0303_ _0304_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_67_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0577_ net27 _0260_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_230_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input129_I la_data_in[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_202_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input94_I la_data_in[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput102 la_data_in[28] net102 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput113 la_data_in[38] net113 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput124 la_data_in[48] net124 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput135 la_data_in[58] net135 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput146 la_data_in[68] net146 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput157 la_data_in[78] net157 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput168 la_data_in[88] net168 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput179 la_data_in[98] net179 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_3911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_57_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_105_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_122_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_220_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput609 net609 la_data_out[86] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0500_ _0202_ _0213_ _0214_ net498 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_214_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_231_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_225_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0662__A4 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0629_ _0232_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_217_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input246_I la_oenb[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input413_I wbs_stb_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1063__A1 _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output632_I net632 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0980_ _0092_ net528 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput417 net417 data_mem_addr[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput428 net428 data_write_data[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput439 net439 data_write_data[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input1_I data_read_data[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1045__A1 _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input196_I la_oenb[113] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input363_I wbs_adr_i[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_11281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input57_I la_data_in[102] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout677 net680 net677 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_130_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout688 net689 net688 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_167_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout699 net42 net699 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1036__A1 net695 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1027__A1 instr_load_addr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0963_ _0224_ _0281_ net473 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_220_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0894_ net495 net172 _0043_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_192_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0561__I0 instr_load_addr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input111_I la_data_in[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input209_I la_oenb[125] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1018__A1 _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_7815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output428_I net428 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0552__I0 _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0983__I _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1009__A1 _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1231_ net404 net671 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1054__I _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1162_ net344 analog_io[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_65_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1093_ _0006_ net706 net681 data_load_addr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XTAP_4091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0946_ _0074_ net513 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0877_ _0035_ net606 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input159_I la_data_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input326_I uP_write_data[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_205_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0773__I0 net456 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0800_ _0410_ net570 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_239_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1082__CLK net681 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0731_ _0352_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_129_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0662_ _0305_ _0310_ _0315_ _0320_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_9581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0593_ net19 _0273_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_8880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0764__I0 net452 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_152_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1214_ net49 net463 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1076_ _0013_ net700 net676 instr_load_addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_59_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0995__A3 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0929_ _0176_ net61 _0064_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_239_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input276_I la_oenb[70] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0798__I _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0755__I0 net633 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput306 la_oenb[98] net306 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput317 uP_dataw_en net317 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_5528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput328 uP_write_data[11] net328 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput339 uP_write_data[7] net339 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_715 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_211_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_726 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_737 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_233_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_748 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xio_interface_759 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_84_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0683__A2 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_246_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output495_I net495 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0746__I0 net629 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0612__S _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0714_ net86 _0345_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_10921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout693_I net440 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0645_ net301 net300 net303 net302 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_10976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0576_ _0263_ _0265_ net635 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_171_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1059_ _0186_ _0153_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input393_I wbs_dat_i[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input87_I la_data_in[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1082__RN net707 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput103 la_data_in[29] net103 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput114 la_data_in[39] net114 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput125 la_data_in[49] net125 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput136 la_data_in[59] net136 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput147 la_data_in[69] net147 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_236_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput158 la_data_in[79] net158 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput169 la_data_in[89] net169 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_107_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_161_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_86_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0967__I0 net693 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_10239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_6571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0607__S _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_143_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_242_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout706_I net710 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0628_ _0293_ net439 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_10795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_214_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0559_ _0187_ net322 _0252_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input141_I la_data_in[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input239_I la_oenb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input406_I wbs_dat_i[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_228_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_241_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output625_I net625 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput418 net418 data_mem_addr[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput429 net429 data_write_data[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_194_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_7080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input189_I la_oenb[107] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input356_I wbs_adr_i[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout678 net679 net678 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_219_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout689 net690 net689 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_21_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1036__A2 _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_221_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_215_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0710__S _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0962_ _0083_ net521 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_207_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0893_ _0044_ net614 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input104_I la_data_in[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0552__I1 net319 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1230_ net403 net670 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_232_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1092_ _0005_ net705 net679 data_load_addr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_228_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0945_ net698 net69 _0070_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0876_ net422 net163 _0033_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_173_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input221_I la_oenb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input319_I uP_instr_mem_addr[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0998__A1 _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0470__I0 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output440_I net691 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput590 net590 la_data_out[69] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0989__A1 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0730_ _0370_ net537 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0661_ _0316_ _0317_ _0318_ _0319_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_155_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_196_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0592_ _0274_ net642 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_8870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1213_ net48 net462 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_242_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1014__B instr_load_addr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1075_ _0012_ net700 net676 instr_load_addr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_91_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0928_ _0048_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_147_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0452__I0 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0859_ net7 net155 _0022_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input171_I la_data_in[90] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input269_I la_oenb[64] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput307 la_oenb[99] net307 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput318 uP_instr_mem_addr[0] net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput329 uP_write_data[12] net329 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input32_I instr[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_716 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xio_interface_727 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_4828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xio_interface_738 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_229_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_749 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_211_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0683__A3 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0691__I0 net409 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output488_I net488 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0713_ _0361_ net529 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_10911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0644_ net296 net295 net299 net298 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_234_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_10966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0575_ _0264_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_136_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1058_ _0137_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input386_I wbs_dat_i[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput104 la_data_in[2] net104 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput115 la_data_in[3] net115 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput126 la_data_in[4] net126 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput137 la_data_in[5] net137 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput148 la_data_in[6] net148 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput159 la_data_in[7] net159 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_241_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_107_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0967__I1 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_225_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0623__S _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0627_ net698 net341 _0289_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_10796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0558_ _0254_ net452 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0489_ net51 net52 _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_189_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input134_I la_data_in[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input301_I la_oenb[93] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0894__I0 net495 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0533__S _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1163__I net355 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0708__S _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0885__I0 net490 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput419 net419 data_mem_addr[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0618__S _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0876__I0 net422 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input251_I la_oenb[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input349_I wbs_adr_i[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout679 net680 net679 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_218_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0867__I0 net418 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output470_I net470 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_237_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_9978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0961_ _0265_ net77 _0080_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0892_ net494 net171 _0043_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_199_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_212_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1018__A3 _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input299_I la_oenb[91] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input62_I la_data_in[107] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_11080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_245_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_196_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1091_ _0004_ net703 net678 data_load_addr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_225_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0944_ _0073_ net512 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0875_ _0034_ net605 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input214_I la_oenb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput580 net580 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput591 net591 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_output433_I net433 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1171__I net375 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0989__A2 _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0660_ net209 net208 net211 net210 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_48_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0591_ net33 _0273_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_9594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_238_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1212_ net47 net461 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1074_ _0008_ net702 net678 instr_load_addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0927_ _0063_ net504 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0601__A1 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0858_ _0024_ net597 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_239_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0789_ _0403_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_170_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input164_I la_data_in[84] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput308 la_oenb[9] net308 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput319 uP_instr_mem_addr[1] net319 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input331_I uP_write_data[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_717 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_22_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_728 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input25_I instr[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xio_interface_739 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_5_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_142_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1166__I net370 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0451__S0 _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0712_ net368 net85 _0358_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0643_ net288 net287 net290 net289 _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_10956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0574_ _0232_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_8690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout679_I net680 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1057_ data_load_addr\[4\] _0150_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input281_I la_oenb[75] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input379_I wbs_dat_i[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput105 la_data_in[30] net105 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput116 la_data_in[40] net116 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput127 la_data_in[50] net127 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput138 la_data_in[60] net138 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput149 la_data_in[70] net149 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0656__A4 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1066__A1 _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_188_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_103_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_224_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0501__C2 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_204_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1057__A1 data_load_addr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_231_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0626_ _0292_ net438 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_10775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0557_ instr_load_addr\[3\] net321 _0252_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_234_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0488_ _0203_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input127_I la_data_in[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1048__A1 _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input92_I la_data_in[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_199_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0523__I data_load_addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0634__S _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout711_I net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_11273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0609_ net35 net333 _0257_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input244_I la_oenb[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0564__I0 _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input411_I wbs_sel_i[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0492__A2 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0544__S _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output463_I net463 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output630_I net630 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1174__I net347 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0555__I0 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_226_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0960_ _0082_ net519 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1085__CLK net685 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0891_ _0027_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_122_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0794__I0 net433 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0546__I0 data_load_addr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input194_I la_oenb[111] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input361_I wbs_adr_i[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_11081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_7818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input55_I la_data_in[100] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_10391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0537__I0 data_load_addr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1169__I net373 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1090_ _0003_ net703 net677 data_load_addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_161_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0943_ net699 net68 _0070_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0874_ net421 net162 _0033_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_239_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_244_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input207_I la_oenb[123] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput570 net570 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_114_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput581 net581 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput592 net592 la_data_out[70] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output426_I net426 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0732__S _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0531__I net694 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0590_ _0237_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_9595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1211_ net46 net460 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1073_ _0163_ net643 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0926_ _0173_ net60 _0059_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0601__A2 _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0857_ net6 net154 _0022_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1094__RN net707 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0441__I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_235_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0788_ _0347_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input157_I la_data_in[78] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput309 uP_data_mem_addr[0] net309 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_233_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xio_interface_718 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_5_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_729 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_217_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input324_I uP_instr_mem_addr[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input18_I instr[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0817__S _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0552__S _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0979__I0 net686 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0451__S1 _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_212_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1182__I net356 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0711_ _0360_ net520 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_10902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0595__A1 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0642_ net292 net291 net294 net293 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_10946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0573_ net26 _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_234_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1056_ data_load_addr\[4\] _0150_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_241_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0909_ _0053_ net621 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0586__A1 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input274_I la_oenb[69] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput106 la_data_in[31] net106 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput117 la_data_in[41] net117 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput128 la_data_in[51] net128 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput139 la_data_in[61] net139 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1066__A2 _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_227_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_107_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_224_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output493_I net493 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_107_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_220_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0577__A1 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1177__I net350 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0501__A1 instr_load_addr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0501__B2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1057__A2 _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout691_I net693 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0625_ net699 net340 _0289_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_10765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0556_ _0253_ net451 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0487_ _0165_ _0167_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1039_ _0137_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1048__A2 _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input391_I wbs_dat_i[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input85_I la_data_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_225_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout704_I net705 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0608_ _0282_ net424 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0539_ data_load_addr\[5\] _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_154_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input237_I la_oenb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input404_I wbs_dat_i[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_243_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output456_I net456 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0555__I1 net320 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1190__I net364 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0890_ _0042_ net612 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0470__S _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0546__I1 net316 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0482__I0 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_8509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input187_I la_oenb[105] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input354_I wbs_adr_i[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_10392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input48_I io_in[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0537__I1 net313 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_230_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0473__I0 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1185__I net359 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_156_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0942_ _0072_ net511 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_220_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0464__I0 _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0873_ _0027_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_103_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_237_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input102_I la_data_in[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_216_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput560 net560 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_161_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput571 net571 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_182_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput582 net582 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput593 net593 la_data_out[71] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output419_I net419 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1210_ net45 net459 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0677__A3 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1072_ net93 net220 _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_1_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0925_ _0062_ net503 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0722__I _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0856_ _0023_ net596 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0787_ _0402_ net564 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_217_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_719 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_211_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input317_I uP_dataw_en vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_107_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0807__I _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_227_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0542__I net694 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0710_ net367 net76 _0358_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0641_ _0300_ net430 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_10936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0572_ _0262_ net634 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_217_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1055_ data_load_addr\[0\] data_load_addr\[1\] data_load_addr\[2\] data_load_addr\[3\]
+ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_213_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_198_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0908_ net485 net178 _0049_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_200_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0830__I0 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0839_ net13 net145 _0431_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input267_I la_oenb[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_227_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput107 la_data_in[32] net107 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput118 la_data_in[42] net118 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput129 la_data_in[52] net129 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input30_I instr[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0510__A2 net695 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_246_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_107_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_161_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_202_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output486_I net486 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_197_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0821__I0 net430 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_180_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1193__I net691 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0738__S _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0812__I0 net426 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_11456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0624_ _0291_ net437 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_9190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout684_I net685 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0555_ _0178_ net320 _0252_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0486_ _0201_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1038_ _0207_ _0168_ _0281_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_179_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input384_I wbs_dat_i[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input78_I la_data_in[121] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0803__I0 net437 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0910__I _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1188__I net362 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0931__S _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0607_ net34 net326 _0257_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_10585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0538_ _0241_ net420 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0469_ _0170_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input132_I la_data_in[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1002__S _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output449_I net449 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput290 la_oenb[83] net290 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_58_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0482__I1 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_11094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input347_I wbs_adr_i[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_180_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0473__I1 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_178_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_210_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0941_ _0198_ net67 _0070_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_222_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0872_ _0032_ net604 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_228_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_177_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input297_I la_oenb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input60_I la_data_in[105] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0463__S0 _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput550 net550 la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput561 net561 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput572 net572 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput583 net583 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_60_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput594 net594 la_data_out[72] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0566__S _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1196__I net692 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0677__A4 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1071_ _0149_ _0161_ _0162_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_198_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0924_ _0164_ net59 _0059_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0855_ net5 net153 _0022_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_200_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0786_ net424 net121 _0392_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1011__A1 _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0445__S0 _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input212_I la_oenb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_146_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output431_I net431 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1069__A1 data_load_addr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0640_ net49 net332 _0264_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_10915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0571_ net25 _0260_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_8660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1054_ _0137_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0907_ _0052_ net620 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_239_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0838_ _0432_ net587 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0769_ net454 net112 _0392_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_46_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input162_I la_data_in[82] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput108 la_data_in[33] net108 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput119 la_data_in[43] net119 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input23_I instr[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_205_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_220_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_224_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_7244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_207_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0623_ net41 net339 _0289_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_10745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0554_ _0244_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_8490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0929__S _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout677_I net680 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0485_ net50 _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1037_ _0116_ _0135_ _0136_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_165_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input377_I wbs_dat_i[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput90 la_data_in[17] net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_217_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0548__I instr_load_addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_11210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_11298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0606_ _0265_ net317 _0223_ _0281_ net440 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_10575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0549__I0 _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0537_ data_load_addr\[4\] net313 _0238_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_234_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0468_ net11 net28 data_load_addr\[4\] _0187_ _0183_ _0179_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input125_I la_data_in[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input90_I la_data_in[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_210_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_194_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_215_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0712__I0 net368 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1199__I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0479__S _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput280 la_oenb[74] net280 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput291 la_oenb[84] net291 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0703__I0 net376 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0482__I2 data_load_addr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0741__I _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_11051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_11073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input242_I la_oenb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output461_I net461 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0933__I0 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0826__I _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0940_ _0071_ net510 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_207_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0871_ net420 net161 _0028_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0924__I0 _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_225_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input192_I la_oenb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0463__S1 _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput540 net540 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_66_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input53_I io_in[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput551 net551 la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput562 net562 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_82_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput573 net573 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_43_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput584 net584 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput595 net595 la_data_out[73] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_219_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0915__I0 net488 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0906__I0 net484 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1070_ _0198_ _0153_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_207_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0923_ _0061_ net502 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1079__RN net702 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0854_ _0425_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_146_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_0785_ _0401_ net563 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_239_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0445__S1 _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0466__I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1199_ net34 net457 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input205_I la_oenb[121] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_142_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output424_I net424 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0570_ _0261_ net627 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_8650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_8661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1053_ _0138_ _0147_ _0148_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_202_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_185_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0906_ net484 net177 _0049_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0837_ net12 net144 _0431_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__0991__A1 _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0768_ _0376_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_85_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0699_ net412 net148 _0353_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input155_I la_data_in[76] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput109 la_data_in[34] net109 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input322_I uP_instr_mem_addr[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input16_I data_read_data[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_107_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output639_I net639 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0498__C2 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_245_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0622_ _0290_ net436 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_10746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0553_ _0251_ net450 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_193_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0484_ _0200_ net496 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_234_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input8_I data_read_data[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1036_ net695 _0114_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input272_I la_oenb[67] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput80 la_data_in[123] net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_116_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput91 la_data_in[18] net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_190_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0919__I _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output491_I net491 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_231_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_11266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0605_ _0170_ net694 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0549__I1 net318 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0536_ _0240_ net419 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0467_ instr_load_addr\[4\] _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_214_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input118_I la_data_in[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1019_ instr_load_addr\[8\] _0121_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_228_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_243_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input83_I la_data_in[126] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput270 la_oenb[65] net270 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_79_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput281 la_oenb[75] net281 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_64_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput292 la_oenb[85] net292 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_111_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout702_I net704 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0482__I3 instr_load_addr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_11041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0519_ _0217_ _0227_ _0228_ net487 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_99_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input235_I la_oenb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input402_I wbs_dat_i[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0458__I0 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0473__I3 instr_load_addr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0630__I0 net697 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output454_I net454 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0870_ _0031_ net603 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_202_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0621__I0 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_205_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0999_ instr_load_addr\[0\] instr_load_addr\[1\] instr_load_addr\[2\] instr_load_addr\[3\]
+ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_238_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input185_I la_oenb[103] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0612__I0 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput530 net530 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput541 net541 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput552 net552 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input352_I wbs_adr_i[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput563 net563 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput574 net574 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput585 net585 la_data_out[64] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input46_I io_in[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput596 net596 la_data_out[74] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_114_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_196_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0773__S _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0922_ _0168_ net58 _0059_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0853_ _0021_ net595 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0784_ net120 _0348_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 data_read_data[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1198_ net440 net448 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_246_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input100_I la_data_in[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output417_I net417 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_207_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1052_ _0182_ _0139_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0905_ _0051_ net619 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0836_ _0425_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_89_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0991__A2 _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0767_ _0391_ net554 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0698_ _0352_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_217_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input148_I la_data_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input315_I uP_data_mem_addr[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_205_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0498__B2 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0621_ net40 net338 _0289_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_10725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0552_ _0250_ net319 _0245_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_8470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0483_ _0198_ _0199_ _0189_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_7780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0489__A1 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_226_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1035_ instr_load_addr\[12\] _0134_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_228_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0961__S _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput70 la_data_in[114] net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_172_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0819_ net429 net136 _0419_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput81 la_data_in[124] net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_46_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput92 la_data_in[19] net92 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_235_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input265_I la_oenb[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0716__A2 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_198_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output484_I net484 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_180_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0845__I _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0604_ _0280_ net633 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_10555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0535_ data_load_addr\[3\] net312 _0238_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_217_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0466_ net38 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_231_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1018_ _0096_ _0119_ _0121_ _0122_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_223_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0691__S _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input382_I wbs_dat_i[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input76_I la_data_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1050__A1 data_load_addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_182_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput260 la_oenb[56] net260 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput271 la_oenb[66] net271 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput282 la_oenb[76] net282 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput293 la_oenb[86] net293 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0575__I _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1041__A1 _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_11042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0518_ _0219_ net48 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0449_ _0172_ net482 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_171_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input130_I la_data_in[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input228_I la_oenb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0485__I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0458__I1 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_221_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1032__A1 net696 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_211_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0998_ _0095_ _0105_ _0106_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1014__A1 _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input178_I la_data_in[97] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput520 net520 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_145_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput531 net531 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput542 net542 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput553 net553 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput564 net564 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput575 net575 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput586 net586 la_data_out[65] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input345_I wbs_adr_i[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput597 net597 la_data_out[75] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_21_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input39_I io_in[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_200_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_8822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0921_ _0060_ net501 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0852_ net4 net152 _0436_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_196_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0783_ _0400_ net562 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_216_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput2 data_read_data[10] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0964__S _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1197_ net693 net447 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_246_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_146_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input295_I la_oenb[88] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0938__I _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_7995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_238_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0760__I0 net450 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1051_ data_load_addr\[3\] _0146_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_228_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0904_ net483 net176 _0049_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0835_ _0430_ net586 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_239_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0766_ net453 net111 _0387_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0959__S _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0697_ _0347_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0751__I0 net631 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1249_ net392 net659 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input210_I la_oenb[126] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input308_I la_oenb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0742__I0 net642 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_201_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0620_ _0232_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_10715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0551_ instr_load_addr\[1\] _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_8460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0482_ net14 net31 data_load_addr\[7\] instr_load_addr\[7\] _0165_ _0167_ _0199_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_7770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0489__A2 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1034_ instr_load_addr\[10\] instr_load_addr\[11\] _0120_ _0126_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_228_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1202__I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0661__A2 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_198_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput60 la_data_in[105] net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_137_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput71 la_data_in[115] net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_0818_ _0420_ net578 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput82 la_data_in[125] net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput93 la_data_in[1] net93 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_217_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0749_ _0381_ net545 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input160_I la_data_in[80] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input258_I la_oenb[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input21_I instr[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0603_ net24 _0233_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_10556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0534_ _0239_ net418 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_8290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0954__I0 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0465_ _0185_ net492 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_224_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1017_ _0198_ _0109_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input375_I wbs_adr_i[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input69_I la_data_in[113] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0945__I0 net698 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1050__A2 _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput250 la_oenb[47] net250 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput261 la_oenb[57] net261 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput272 la_oenb[67] net272 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput283 la_oenb[77] net283 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput294 la_oenb[87] net294 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0792__S _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1041__A2 _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_11032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_11043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0967__S _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0517_ net6 _0223_ _0224_ net23 _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_154_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0448_ _0164_ _0169_ _0171_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input123_I la_data_in[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0458__I2 _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1032__A2 _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_237_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1210__I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0997_ _0182_ _0099_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput510 net510 la_data_out[110] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput521 net521 la_data_out[120] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput532 net532 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput543 net543 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput554 net554 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_236_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput565 net565 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput576 net576 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput587 net587 la_data_out[66] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_113_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput598 net598 la_data_out[76] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_60_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input240_I la_oenb[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input338_I uP_write_data[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1005__A2 instr_load_addr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_9579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0920_ _0166_ net57 _0059_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0851_ _0439_ net594 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0782_ net119 _0396_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_100_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_237_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1205__I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput3 data_read_data[11] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1196_ net692 net446 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0994__A1 _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input190_I la_oenb[108] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input288_I la_oenb[81] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input51_I io_in[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_240_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0985__A1 _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_9387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1050_ data_load_addr\[0\] _0235_ _0177_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_111_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0864__I _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0903_ _0050_ net618 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0834_ net11 net143 _0426_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_200_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0765_ _0390_ net553 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0696_ _0351_ net580 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0975__S _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1248_ net391 net658 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1179_ net352 analog_io[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_38_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input203_I la_oenb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input99_I la_data_in[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output422_I net422 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_204_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0550_ _0249_ net449 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_234_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0481_ net41 _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_234_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_238_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1033_ _0116_ _0132_ _0133_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_207_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput50 io_in[32] net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_176_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput61 la_data_in[106] net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_0817_ net428 net135 _0419_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput72 la_data_in[116] net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_50_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput83 la_data_in[126] net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_239_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput94 la_data_in[20] net94 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_157_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0748_ net630 net102 _0377_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0679_ net235 net234 net237 net236 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_22_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input153_I la_data_in[74] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input320_I uP_instr_mem_addr[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input14_I data_read_data[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_199_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_7012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output637_I net637 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput410 wbs_sel_i[1] net410 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0479__I0 _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0602_ _0279_ net632 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_10535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0533_ _0177_ net311 _0238_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_234_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0464_ _0182_ _0184_ _0171_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_7590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input6_I data_read_data[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1213__I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1016_ _0120_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_165_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input270_I la_oenb[65] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input368_I wbs_adr_i[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0962__I _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1050__A3 _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput240 la_oenb[38] net240 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput251 la_oenb[48] net251 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput262 la_oenb[58] net262 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_79_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput273 la_oenb[68] net273 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput284 la_oenb[78] net284 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput295 la_oenb[88] net295 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1208__I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0516_ _0217_ _0225_ _0226_ net486 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0447_ _0170_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_3_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input116_I la_data_in[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0458__I3 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_9706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input81_I la_data_in[124] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout700_I net702 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0996_ instr_load_addr\[3\] _0104_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_192_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput500 net500 la_data_out[101] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_138_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput511 net511 la_data_out[111] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput522 net522 la_data_out[121] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput533 net533 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_216_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput544 net544 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput555 net555 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput566 net566 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_233_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput577 net577 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput588 net588 la_data_out[67] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_5_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput599 net599 la_data_out[77] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input233_I la_oenb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input400_I wbs_dat_i[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output452_I net452 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_8868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0850_ net3 net151 _0436_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0781_ _0399_ net561 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0507__A2 net696 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_155_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 data_read_data[12] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1195_ net692 net445 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_209_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0979_ net686 net84 _0344_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_238_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input183_I la_oenb[101] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input350_I wbs_adr_i[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input44_I io_in[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0985__A2 _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_240_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0902_ net498 net175 _0049_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_19_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0833_ _0429_ net585 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0764_ net452 net110 _0387_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout698_I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0695_ net411 net137 _0348_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1216__I net690 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1247_ net390 net657 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1178_ net351 analog_io[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_181_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_59_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input398_I wbs_dat_i[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0965__I _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output415_I net686 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_245_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_201_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0480_ _0197_ net495 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_234_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1032_ net696 _0114_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_235_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0661__A4 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1071__A1 _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput40 io_in[22] net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0816_ _0403_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput51 io_in[33] net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput62 la_data_in[107] net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput73 la_data_in[117] net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_89_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput84 la_data_in[127] net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_196_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput95 la_data_in[21] net95 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0747_ _0380_ net544 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0678_ net239 net238 net241 net240 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_233_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input146_I la_data_in[68] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_211_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input313_I uP_data_mem_addr[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1062__A1 _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput400 wbs_dat_i[30] net400 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput411 wbs_sel_i[2] net411 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_207_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_207_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1053__A1 _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0601_ net23 _0233_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_10525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0532_ _0237_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_8270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0463_ net10 net27 data_load_addr\[3\] instr_load_addr\[3\] _0183_ _0179_ _0184_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_7580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1015_ instr_load_addr\[6\] instr_load_addr\[7\] _0107_ _0112_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_143_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1044__A1 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0478__S0 _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input263_I la_oenb[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output482_I net482 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1035__A1 instr_load_addr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_216_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput230 la_oenb[29] net230 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_40_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput241 la_oenb[39] net241 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput252 la_oenb[49] net252 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput263 la_oenb[59] net263 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput274 la_oenb[69] net274 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput285 la_oenb[79] net285 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_236_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput296 la_oenb[89] net296 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1026__A1 _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_11001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_11045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0515_ _0219_ net47 _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_fanout680_I net684 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0446_ net50 _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_234_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1224__I net711 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input109_I la_data_in[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1017__A1 _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input380_I wbs_dat_i[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input74_I la_data_in[118] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1008__A1 _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0790__I0 net431 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0995_ instr_load_addr\[0\] _0250_ _0178_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_14_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput501 net501 la_data_out[102] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput512 net512 la_data_out[112] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_157_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput523 net523 la_data_out[122] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_218_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput534 net534 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput545 net545 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput556 net556 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput567 net567 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_86_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput578 net578 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput589 net589 la_data_out[68] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_29_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input226_I la_oenb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0533__I0 _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_9526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0968__I _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0780_ net118 _0396_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1039__I _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput5 data_read_data[13] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1194_ net692 net444 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0978_ _0091_ net415 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1081__CLK net681 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input176_I la_data_in[95] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0788__I _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_190_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input343_I wb_rst_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input37_I io_in[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0682__A2 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0698__I _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_215_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0901_ _0048_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_203_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0832_ net10 net142 _0426_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0763_ _0389_ net552 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0694_ _0350_ net569 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0736__I0 net640 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1246_ net389 net656 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_246_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1177_ net350 analog_io[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input293_I la_oenb[86] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0975__I0 net342 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1081__RN net707 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0727__I0 net636 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0591__A1 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_8496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1031_ instr_load_addr\[11\] _0131_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0646__A2 _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_185_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0891__I _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput30 instr[6] net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput41 io_in[23] net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_201_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0815_ _0418_ net577 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput52 io_in[34] net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_239_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput63 la_data_in[108] net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput74 la_data_in[118] net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_176_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput85 la_data_in[12] net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_0746_ net629 net101 _0377_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput96 la_data_in[22] net96 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_85_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0957__I0 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0582__A1 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0677_ _0332_ _0333_ _0334_ _0335_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_26_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input139_I la_data_in[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1229_ net402 net669 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input306_I la_oenb[98] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1062__A2 _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0948__I0 net697 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_231_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput401 wbs_dat_i[31] net401 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput412 wbs_sel_i[3] net412 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_196_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_236_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_199_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_240_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0600_ _0278_ _0265_ net631 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_138_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0939__I0 _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0531_ net694 _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_8260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0462_ _0165_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_7570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1014_ _0195_ _0113_ instr_load_addr\[7\] _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_1_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1044__A2 _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_236_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0729_ net637 net94 _0366_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_235_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input256_I la_oenb[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_228_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output642_I net642 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput220 la_oenb[1] net220 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput231 la_oenb[2] net231 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput242 la_oenb[3] net242 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_20_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput253 la_oenb[4] net253 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput264 la_oenb[5] net264 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput275 la_oenb[6] net275 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput286 la_oenb[7] net286 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput297 la_oenb[8] net297 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_223_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_220_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_11068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0514_ net5 _0223_ _0224_ net22 _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_8090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0445_ net1 net18 data_load_addr\[0\] instr_load_addr\[0\] _0166_ _0168_ _0169_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_80_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1017__A2 _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input373_I wbs_adr_i[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input67_I la_data_in[111] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_210_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1008__A2 _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_237_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_159_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0994_ _0095_ _0102_ _0103_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput502 net502 la_data_out[103] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput513 net513 la_data_out[113] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_216_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput524 net524 la_data_out[123] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput535 net535 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput546 net546 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_236_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput557 net557 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput568 net568 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput579 net579 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_87_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__0533__I1 net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input121_I la_data_in[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input219_I la_oenb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0997__A1 _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output438_I net438 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0984__I _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_210_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 data_read_data[14] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_5080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1193_ net691 net443 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1004__B instr_load_addr\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0977_ net54 net342 _0264_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_238_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0451__I0 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input169_I la_data_in[89] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input336_I uP_write_data[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_7933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_8689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_0900_ _0424_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0831_ _0428_ net584 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0762_ net451 net109 _0387_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_196_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0693_ net410 net126 _0348_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_9891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1245_ net387 net654 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_228_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1176_ net349 analog_io[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input286_I la_oenb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_7207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_210_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_10708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1030_ instr_load_addr\[10\] _0121_ _0126_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_169_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput20 instr[11] net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput31 instr[7] net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_0814_ net427 net134 _0414_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_190_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput42 io_in[24] net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput53 io_in[36] net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_217_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput64 la_data_in[109] net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput75 la_data_in[119] net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_50_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0745_ _0379_ net543 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput86 la_data_in[13] net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput97 la_data_in[23] net97 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_67_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0676_ net266 net265 net268 net267 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_63_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1228_ net399 net666 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input201_I la_oenb[118] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input97_I la_data_in[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_7037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput402 wbs_dat_i[3] net402 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput413 wbs_stb_i net413 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output420_I net420 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_145_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0636__I0 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_156_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0530_ _0236_ net417 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_8250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0461_ net37 _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_7560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1013_ _0116_ _0117_ _0118_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_228_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0627__I0 net698 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0728_ _0369_ net536 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_232_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0659_ net205 net204 net207 net206 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_154_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input151_I la_data_in[72] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input249_I la_oenb[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input12_I data_read_data[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0618__I0 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output468_I net468 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_159_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_235_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output635_I net635 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput210 la_oenb[126] net210 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput221 la_oenb[20] net221 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_6188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput232 la_oenb[30] net232 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput243 la_oenb[40] net243 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput254 la_oenb[50] net254 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput265 la_oenb[60] net265 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput276 la_oenb[70] net276 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput287 la_oenb[80] net287 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput298 la_oenb[90] net298 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0857__I0 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_207_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0609__I0 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_103_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1058__I _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_11047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0513_ _0208_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_8080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0444_ _0167_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_7390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input4_I data_read_data[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0848__I0 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input199_I la_oenb[116] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input366_I wbs_adr_i[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0839__I0 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_202_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_226_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0993_ _0176_ _0099_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0621__S _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput503 net503 la_data_out[104] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput514 net514 la_data_out[114] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_246_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput525 net525 la_data_out[124] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_114_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput536 net536 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_237_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput547 net547 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_218_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput558 net558 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput569 net569 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input114_I la_data_in[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0997__A2 _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput7 data_read_data[15] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1192_ net691 net442 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0616__S _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0976_ _0090_ net527 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0451__I1 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input231_I la_oenb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input329_I uP_write_data[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_227_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0682__A4 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0526__S _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output450_I net450 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_8657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0830_ net9 net141 _0426_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0761_ _0388_ net551 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0692_ _0349_ net558 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_237_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1244_ net386 net653 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1175_ net348 analog_io[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_59_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0959_ net49 net75 _0080_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input181_I la_data_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input279_I la_oenb[73] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input42_I io_in[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output498_I net498 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_199_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_211_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_7775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1056__A1 data_load_addr\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput10 data_read_data[3] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_238_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput21 instr[12] net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_204_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0813_ _0417_ net576 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput32 instr[8] net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput43 io_in[25] net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput54 io_in[37] net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_176_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput65 la_data_in[10] net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_0744_ net628 net100 _0377_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput76 la_data_in[11] net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_89_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput87 la_data_in[14] net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_196_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput98 la_data_in[24] net98 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout696_I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_154_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0675_ net261 net260 net263 net262 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_48_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1227_ net388 net655 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1089_ _0002_ net701 net677 data_load_addr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_33_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1047__A1 _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input396_I wbs_dat_i[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput403 wbs_dat_i[4] net403 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_66_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput414 wbs_we_i net414 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_189_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_220_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_142_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_10528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0460_ _0181_ net490 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_171_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1012_ _0194_ _0099_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1029__A1 _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout709_I net710 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0727_ net636 net92 _0366_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_200_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0658_ net196 net195 net198 net197 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0589_ _0272_ net641 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input144_I la_data_in[66] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input311_I uP_data_mem_addr[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input409_I wbs_sel_i[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output628_I net628 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1164__I net366 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput200 la_oenb[117] net200 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput211 la_oenb[127] net211 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_42_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput222 la_oenb[21] net222 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput233 la_oenb[31] net233 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput244 la_oenb[41] net244 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput255 la_oenb[51] net255 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput266 la_oenb[61] net266 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput277 la_oenb[71] net277 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput288 la_oenb[81] net288 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput299 la_oenb[91] net299 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0512_ _0205_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_8070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0443_ net52 _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_218_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1084__CLK net685 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input261_I la_oenb[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input359_I wbs_adr_i[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_154_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0529__S _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output480_I net480 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0992_ _0178_ _0101_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_203_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_10111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput504 net504 la_data_out[105] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput515 net515 la_data_out[115] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput526 net526 la_data_out[125] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput537 net537 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput548 net548 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput559 net559 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_233_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0766__I0 net453 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input107_I la_data_in[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input72_I la_data_in[116] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_8817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0757__I0 net449 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0748__I0 net630 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1191_ net691 net441 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput8 data_read_data[1] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_228_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0920__I0 _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0975_ net342 net83 _0344_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__0632__S _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0600__A2 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0451__I2 data_load_addr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1093__RN net706 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input224_I la_oenb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0667__A2 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0911__I0 net486 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_216_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1172__I net345 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0902__I0 net498 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_245_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_163_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0452__S _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0760_ net450 net108 _0387_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_183_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0969__I0 net317 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0691_ net409 net115 _0348_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_9871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1243_ net385 net652 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1174_ net347 analog_io[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0627__S _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0958_ _0081_ net518 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0889_ net493 net169 _0038_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_7209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input174_I la_data_in[93] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input341_I uP_write_data[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input35_I io_in[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0537__S _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1167__I net371 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0500__A1 _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1056__A2 _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput11 data_read_data[4] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_0812_ net426 net133 _0414_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput22 instr[13] net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput33 instr[9] net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput44 io_in[26] net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_201_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput55 la_data_in[100] net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput66 la_data_in[110] net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_0743_ _0378_ net542 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput77 la_data_in[120] net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_217_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_217_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput88 la_data_in[15] net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput99 la_data_in[25] net99 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_171_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0674_ net252 net251 net255 net254 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout689_I net690 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_230_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1226_ net377 net644 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1088_ _0001_ net701 net676 data_load_addr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input291_I la_oenb[84] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input389_I wbs_dat_i[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput404 wbs_dat_i[5] net404 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0494__C2 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_231_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1038__A2 _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1011_ _0195_ _0113_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_235_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0640__S _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0726_ _0368_ net535 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_154_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0657_ net200 net199 net202 net201 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_170_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0588_ net32 _0268_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_230_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input137_I la_data_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1209_ net44 net458 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input304_I la_oenb[96] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput201 la_oenb[118] net201 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_81_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput212 la_oenb[12] net212 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput223 la_oenb[22] net223 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_194_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput234 la_oenb[32] net234 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput245 la_oenb[42] net245 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_40_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput256 la_oenb[52] net256 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_44_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput267 la_oenb[62] net267 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput278 la_oenb[72] net278 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput289 la_oenb[82] net289 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1180__I net353 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0524__I net694 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_158_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_11038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0511_ _0217_ _0221_ _0222_ net485 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_8060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0442_ _0165_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_7370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0709_ _0359_ net509 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input254_I la_oenb[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output473_I net690 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output640_I net640 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1175__I net348 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0991_ _0248_ _0250_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_220_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0463__I0 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput505 net505 la_data_out[106] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput516 net516 la_data_out[116] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_218_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput527 net527 la_data_out[126] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput538 net538 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput549 net549 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_149_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input371_I wbs_adr_i[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_8818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_8829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input65_I la_data_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_11380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout710 net711 net710 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0693__I0 net410 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0445__I0 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1190_ net364 analog_io[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput9 data_read_data[2] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0974_ _0089_ net526 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0451__I3 instr_load_addr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input217_I la_oenb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_196_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0823__S _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_221_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output436_I net436 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_145_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0532__I _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0690_ _0347_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_9861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1242_ net384 net651 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1173_ net346 analog_io[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_2_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0707__I _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0957_ net48 net74 _0080_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0888_ _0041_ net611 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input167_I la_data_in[87] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input334_I uP_write_data[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input28_I instr[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0896__I0 net496 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_244_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0576__A2 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_7755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1183__I net357 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0887__I0 net492 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0811_ _0416_ net575 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput12 data_read_data[5] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput23 instr[14] net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput34 io_in[16] net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput45 io_in[27] net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0742_ net642 net99 _0377_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_217_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput56 la_data_in[101] net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput67 la_data_in[111] net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput78 la_data_in[121] net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_176_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput89 la_data_in[16] net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0673_ net257 net256 net259 net258 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_9691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1225_ net53 net626 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__0638__S _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0878__I0 net423 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1087_ _0000_ net700 net676 data_load_addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input284_I la_oenb[78] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0900__I _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput405 wbs_dat_i[6] net405 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0869__I0 net419 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0494__B2 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_224_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1038__A3 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_246_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_237_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1178__I net351 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_11209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1010_ _0094_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0725_ net635 net91 _0366_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_171_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0656_ _0311_ _0312_ _0313_ _0314_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_83_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0587_ _0271_ net640 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1208_ net43 net472 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input95_I la_data_in[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput202 la_oenb[119] net202 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_1_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput213 la_oenb[13] net213 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput224 la_oenb[23] net224 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput235 la_oenb[33] net235 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput246 la_oenb[43] net246 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_79_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput257 la_oenb[53] net257 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput268 la_oenb[63] net268 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput279 la_oenb[73] net279 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_207_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_199_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_103_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_194_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0510_ _0219_ net695 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0441_ net51 _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_7360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0450__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_239_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0708_ net365 net65 _0358_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_10872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0639_ _0299_ net429 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_232_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input247_I la_oenb[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_225_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input414_I wbs_we_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input10_I data_read_data[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output633_I net633 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1191__I net691 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_209_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0736__S _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0990_ _0095_ _0098_ _0100_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_203_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0463__I1 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput506 net506 la_data_out[107] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput517 net517 la_data_out[117] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput528 net528 la_data_out[127] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput539 net539 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_237_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I data_read_data[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0603__A1 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input197_I la_oenb[114] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input364_I wbs_adr_i[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_11381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input58_I la_data_in[103] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout700 net702 net700 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_10691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout711 net343 net711 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_243_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_230_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0445__I1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1186__I net360 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0973_ net54 net82 _0085_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input112_I la_data_in[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output429_I net429 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_189_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1068__A1 _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_204_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_208_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1241_ net383 net650 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1172_ net345 analog_io[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1059__A1 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0956_ _0069_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_179_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0887_ net492 net168 _0038_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input327_I uP_write_data[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0810_ net425 net132 _0414_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput13 data_read_data[6] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_223_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput24 instr[15] net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_204_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput35 io_in[17] net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput46 io_in[28] net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
X_0741_ _0376_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput57 la_data_in[102] net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_156_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput68 la_data_in[112] net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput79 la_data_in[122] net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_158_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0672_ _0327_ _0328_ _0329_ _0330_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_67_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_211_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1224_ net711 net625 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1086_ _0011_ net708 net685 instr_load_addr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0939_ _0194_ net66 _0070_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input277_I la_oenb[71] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input40_I io_in[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0566__I0 instr_load_addr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput406 wbs_dat_i[7] net406 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_66_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0564__S _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_220_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output496_I net496 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_145_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_181_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_8210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1194__I net692 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_8265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0557__I0 instr_load_addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0474__S _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0724_ _0367_ net534 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0796__I0 net434 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout694_I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0655_ net191 net190 net194 net193 _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0586_ net31 _0268_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1207_ net42 net471 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0720__I0 net627 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1069_ data_load_addr\[7\] _0160_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_165_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input394_I wbs_dat_i[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input88_I la_data_in[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_235_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput203 la_oenb[11] net203 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput214 la_oenb[14] net214 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_44_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput225 la_oenb[24] net225 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput236 la_oenb[34] net236 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput247 la_oenb[44] net247 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput258 la_oenb[54] net258 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput269 la_oenb[64] net269 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_232_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1189__I net363 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_240_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0440_ net34 _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_8095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_7394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0950__I0 net696 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout707_I net709 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0731__I _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0769__I0 net454 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0707_ _0352_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_10851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0638_ net48 net331 _0264_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_10895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0569_ net18 _0260_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input142_I la_data_in[64] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0941__I0 _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input407_I wbs_dat_i[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_237_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output626_I net626 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0816__I _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0463__I2 data_load_addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0551__I instr_load_addr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput507 net507 la_data_out[108] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput518 net518 la_data_out[118] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_29_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput529 net529 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_5_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_214_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0603__A2 _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_203_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0461__I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_8809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input357_I wbs_adr_i[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout701 net702 net701 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0445__I2 data_load_addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_196_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_229_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0972_ _0088_ net525 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0597__A1 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1078__RN net705 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input105_I la_data_in[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0588__A1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input70_I la_data_in[114] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_226_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_230_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_180_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0579__A1 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1197__I net693 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1240_ net382 net649 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1171_ net375 analog_io[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_20_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0503__A1 _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_237_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1059__A2 _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0955_ _0079_ net517 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0886_ _0040_ net610 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0990__A1 _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input222_I la_oenb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_235_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_202_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 data_read_data[7] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput25 instr[1] net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_239_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput36 io_in[18] net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_0740_ _0347_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput47 io_in[29] net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_141_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput58 la_data_in[103] net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput69 la_data_in[113] net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_217_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0671_ net308 net297 net203 net192 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_9671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_196_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1223_ net17 net491 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0935__S _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1085_ _0010_ net708 net685 instr_load_addr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_181_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0938_ _0069_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_198_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0869_ net419 net160 _0028_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0963__A1 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input172_I la_data_in[91] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput407 wbs_dat_i[8] net407 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input33_I instr[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output489_I net489 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_7521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0557__I1 net321 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0723_ net634 net90 _0366_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0654_ net187 net186 net189 net188 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_28_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0585_ _0270_ net639 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1206_ net41 net470 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1068_ _0242_ data_load_addr\[6\] _0151_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_55_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input387_I wbs_dat_i[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput204 la_oenb[120] net204 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput215 la_oenb[15] net215 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_24_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput226 la_oenb[25] net226 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_216_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput237 la_oenb[35] net237 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput248 la_oenb[45] net248 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_40_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput259 la_oenb[55] net259 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1077__CLK net677 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0706_ _0357_ net624 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0637_ _0298_ net428 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_10885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0568_ _0237_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0499_ _0211_ net698 _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input135_I la_data_in[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input302_I la_oenb[94] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0606__B1 _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output521_I net521 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0448__I0 _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0463__I3 instr_load_addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_196_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput508 net508 la_data_out[109] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput519 net519 la_data_out[119] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_225_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input252_I la_oenb[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout702 net704 net702 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0445__I3 instr_load_addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__0850__I0 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_178_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0827__I _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0971_ net711 net81 _0085_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0841__I0 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0521__A2 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_227_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0472__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0832__I0 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input63_I la_data_in[108] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_11180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0823__I0 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_196_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1170_ net374 analog_io[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_94_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0954_ net47 net73 _0075_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_242_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0814__I0 net427 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0885_ net490 net167 _0038_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input215_I la_oenb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0805__I0 net438 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0981__A2 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_8448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output434_I net434 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0497__A1 _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput15 data_read_data[8] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput26 instr[2] net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput37 io_in[19] net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_201_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput48 io_in[30] net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput59 la_data_in[104] net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_0670_ net213 net212 net215 net214 _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_9650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1222_ net688 net481 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1084_ _0009_ net708 net685 instr_load_addr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_228_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0937_ _0424_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0750__I _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0868_ _0030_ net601 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__0963__A2 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0799_ net435 net127 _0409_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_6309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input165_I la_data_in[85] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_217_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput408 wbs_dat_i[9] net408 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input332_I uP_write_data[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input26_I instr[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_151_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_181_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_8212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_234_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0771__S _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0570__I _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0722_ _0352_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0653_ net305 net304 net307 net306 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_63_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0584_ net30 _0268_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_170_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1205_ net40 net469 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1067_ _0149_ _0158_ _0159_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_198_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input282_I la_oenb[76] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput205 la_oenb[121] net205 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput216 la_oenb[16] net216 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput227 la_oenb[26] net227 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput238 la_oenb[36] net238 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput249 la_oenb[46] net249 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_79_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_235_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_8075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0705_ net413 net181 _0353_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_11576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0636_ net47 net330 _0294_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_10886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0567_ _0259_ net456 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0498_ instr_load_addr\[9\] _0204_ _0206_ net16 _0209_ net33 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input128_I la_data_in[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0606__A1 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0606__B2 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input93_I la_data_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1031__A1 instr_load_addr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput509 net509 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_5_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_10138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_6492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1013__A1 _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_11351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout703 net704 net703 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_63_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0619_ _0288_ net435 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_193_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input245_I la_oenb[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_210_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input412_I wbs_sel_i[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_208_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output464_I net464 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1004__A1 _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_172_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output631_I net631 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0970_ _0087_ net524 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_233_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input195_I la_oenb[112] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_238_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_11170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input362_I wbs_adr_i[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_11181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_11192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input56_I la_data_in[101] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0928__I _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_204_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_243_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_243_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_228_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0573__I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0953_ _0078_ net516 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0884_ _0039_ net609 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input110_I la_data_in[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input208_I la_oenb[124] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_181_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_203_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput670 net670 wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_153_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output427_I net427 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput16 data_read_data[9] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput27 instr[3] net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_196_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput38 io_in[20] net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput49 io_in[31] net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_217_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_217_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0769__S _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0568__I _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1221_ net687 net480 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0732__I0 net638 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1083_ _0020_ net707 net682 instr_load_addr\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_185_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0936_ _0068_ net508 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0799__I0 net435 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_179_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0867_ net418 net158 _0028_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0798_ _0403_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input158_I la_data_in[79] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput409 wbs_sel_i[0] net409 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__0971__I0 net711 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input325_I uP_instr_mem_addr[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0723__I0 net634 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input19_I instr[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_246_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0651__A2 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_8202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0721_ _0365_ net533 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0652_ net183 net182 net185 net184 _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_9481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0583_ _0269_ net638 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_8780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_214_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1204_ net39 net468 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0705__I0 net413 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1066_ _0194_ _0153_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_228_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_202_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0919_ _0048_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input275_I la_oenb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput206 la_oenb[122] net206 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput217 la_oenb[17] net217 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput228 la_oenb[27] net228 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput239 la_oenb[37] net239 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_231_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_246_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_181_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output494_I net494 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_184_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0935__I0 _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0581__I _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0704_ _0356_ net613 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0635_ _0297_ net427 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout692_I net693 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0566_ instr_load_addr\[7\] net325 _0257_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0926__I0 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0957__S _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0497_ _0202_ _0210_ _0212_ net497 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_6_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1049_ _0138_ _0144_ _0145_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0606__A2 net317 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0491__I net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input392_I wbs_dat_i[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input86_I la_data_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0917__I0 _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1022__A2 _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0908__I0 net485 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout705_I net706 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_176_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1200__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_148_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_11385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0618_ net39 net337 _0284_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_10695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout704 net705 net704 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_150_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0549_ _0248_ net318 _0245_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input140_I la_data_in[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input238_I la_oenb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_215_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input405_I wbs_dat_i[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1004__A2 _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_218_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0993__A1 _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input188_I la_oenb[106] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input355_I wbs_adr_i[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_236_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input49_I io_in[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_93_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_243_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_243_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_210_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_194_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_9822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0854__I _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0790__S _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0952_ net695 net72 _0075_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0883_ net489 net166 _0038_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_220_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_233_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_233_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_229_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input103_I la_data_in[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput660 net660 wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput671 net671 wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput17 hlt net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xinput28 instr[4] net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_204_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput39 io_in[21] net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1220_ net687 net479 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1082_ _0019_ net707 net681 instr_load_addr\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_4_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0935_ _0191_ net64 _0064_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_239_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0866_ _0029_ net600 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_220_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0797_ _0408_ net568 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0759__I _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0695__S _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input220_I la_oenb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input318_I uP_instr_mem_addr[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_168_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_205_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_180_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput490 net490 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_160_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0478__I0 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0720_ net627 net89 _0358_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_239_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0651_ _0306_ _0307_ _0308_ _0309_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0582_ net29 _0268_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_8770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1203_ net38 net467 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_238_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1065_ data_load_addr\[6\] _0157_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_230_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1203__I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0918_ _0058_ net500 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_239_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0849_ _0438_ net593 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input170_I la_data_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input268_I la_oenb[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_157_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput207 la_oenb[123] net207 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_79_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput218 la_oenb[18] net218 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_44_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput229 la_oenb[28] net229 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input31_I instr[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_224_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_246_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0880__I0 net482 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output487_I net487 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0632__I0 net696 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_8000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0699__I0 net412 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0871__I0 net420 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0623__I0 net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0703_ net376 net170 _0353_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_11556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0634_ net695 net329 _0294_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_10866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0565_ _0258_ net455 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_fanout685_I net686 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0496_ _0211_ net699 _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_234_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_241_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0973__S _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1048_ _0176_ _0139_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_241_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input385_I wbs_dat_i[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0614__I0 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input79_I la_data_in[122] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0947__I _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_194_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_6461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1090__CLK net677 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_242_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_10630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0617_ _0287_ net434 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_217_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout705 net706 net705 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_10696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0548_ instr_load_addr\[0\] _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0479_ _0194_ _0196_ _0189_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input133_I la_data_in[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input300_I la_oenb[92] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0515__A2 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_236_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput390 wbs_dat_i[21] net390 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_40_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_244_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1211__I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_211_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0817__I0 net428 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0993__A2 _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input250_I la_oenb[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input348_I wbs_adr_i[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_3_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_3_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_243_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0808__I0 net439 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_204_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_194_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0672__A1 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0951_ _0077_ net515 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0882_ _0027_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_51_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1206__I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input298_I la_oenb[90] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input61_I la_data_in[106] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0718__A2 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput650 net650 wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_236_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput661 net661 wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_82_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput672 net672 wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_156_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_240_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0690__I _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput18 instr[0] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput29 instr[5] net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_32_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1081_ _0018_ net707 net681 instr_load_addr\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0934_ _0067_ net507 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1070__A1 _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0865_ net417 net157 _0028_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_200_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0796_ net434 net125 _0404_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_233_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0775__I _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_183_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input213_I la_oenb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_209_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1061__A1 _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput480 net480 instrw_en_8bit[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_216_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput491 net491 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output432_I net432 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0478__I1 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1052__A1 _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0650_ net283 net282 net285 net284 _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_9461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0581_ _0237_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_8760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0796__S _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1202_ net37 net466 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_230_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1064_ _0242_ _0151_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1043__A1 _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0917_ _0202_ net56 _0054_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0848_ net2 net150 _0436_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0779_ _0398_ net560 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input163_I la_data_in[83] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput208 la_oenb[124] net208 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput219 la_oenb[19] net219 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA_input330_I uP_write_data[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input24_I instr[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_244_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_205_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1034__A1 instr_load_addr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0468__S0 _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1025__A1 net698 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0702_ _0355_ net602 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_11546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0633_ _0296_ net426 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_10845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0564_ _0195_ net324 _0257_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_8590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0495_ net50 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1214__I net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1047_ _0177_ _0143_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_241_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input280_I la_oenb[74] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_175_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input378_I wbs_dat_i[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0873__I _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1209__I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_11387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0616_ net38 net336 _0284_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_10675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_10697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0509__C2 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout706 net710 net706 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_214_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0547_ _0247_ net423 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_230_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0478_ net13 net30 data_load_addr\[6\] _0195_ _0183_ _0167_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input126_I la_data_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input91_I la_data_in[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0771__I0 net455 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0762__I0 net451 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput380 wbs_dat_i[12] net380 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_75_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput391 wbs_dat_i[22] net391 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_212_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_229_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_203_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout710_I net711 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0979__S _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_11173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input243_I la_oenb[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0753__I0 net632 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input410_I wbs_sel_i[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_230_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_243_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_196_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output462_I net462 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1080__CLK net681 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_219_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_9857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0744__I0 net628 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_150_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0950_ net696 net71 _0075_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0881_ _0037_ net608 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_242_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input193_I la_oenb[110] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_197_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input360_I wbs_adr_i[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput640 net640 uP_instr[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_160_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input54_I io_in[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput651 net651 wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput662 net662 wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput673 net673 wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1080__RN net705 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_210_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput19 instr[10] net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_8942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1080_ _0017_ net705 net681 instr_load_addr\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_130_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0933_ _0186_ net63 _0064_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1070__A2 _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0864_ _0027_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_89_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0795_ _0407_ net567 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0708__I0 net365 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input206_I la_oenb[122] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_205_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput470 net470 instr_write_data[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_156_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput481 net481 instrw_en_8bit[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput492 net492 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0966__I _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output425_I net425 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1052__A2 _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0580_ _0267_ net637 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_9495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1201_ net36 net465 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1063_ _0149_ _0155_ _0156_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1043__A2 _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0916_ _0057_ net499 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0847_ _0437_ net592 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_239_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0929__I0 _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0778_ net117 _0396_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_44_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input156_I la_data_in[77] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput209 la_oenb[125] net209 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_211_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input323_I uP_instr_mem_addr[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input17_I hlt vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_103_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1034__A2 instr_load_addr\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0468__S1 _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_194_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1025__A2 _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_184_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0701_ net414 net159 _0353_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_11536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_10802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0632_ net696 net328 _0294_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_10835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0563_ _0244_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_8580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0494_ instr_load_addr\[8\] _0204_ _0206_ net15 _0209_ net32 _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XTAP_7890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I data_read_data[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_230_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1046_ _0231_ _0235_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_200_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input273_I la_oenb[68] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_162_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_213_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output492_I net492 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_205_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_245_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0615_ _0286_ net433 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_236_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0509__A1 instr_load_addr\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0509__B2 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout707 net709 net707 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0546_ data_load_addr\[7\] net316 _0245_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_234_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1225__I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0477_ instr_load_addr\[6\] _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_214_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input119_I la_data_in[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1029_ _0116_ _0129_ _0130_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_241_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0996__A1 instr_load_addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input390_I wbs_dat_i[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input84_I la_data_in[127] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_202_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_246_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0987__A1 _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_164_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput370 wbs_adr_i[4] net370 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput381 wbs_dat_i[13] net381 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_20_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput392 wbs_dat_i[23] net392 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout703_I net704 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_242_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_11174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0529_ _0235_ net310 _0233_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input236_I la_oenb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input403_I wbs_dat_i[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_243_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_243_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output455_I net455 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_246_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0880_ net482 net165 _0033_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_196_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input186_I la_oenb[104] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0789__I _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput630 net630 uP_instr[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_172_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput641 net641 uP_instr[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput652 net652 wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input353_I wbs_adr_i[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput663 net663 wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput674 net674 wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input47_I io_in[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_214_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_211_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_8998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0932_ _0066_ net506 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0863_ _0424_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_204_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0794_ net433 net124 _0404_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_192_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_237_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_246_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_224_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input101_I la_data_in[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__0892__I0 net494 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput460 net460 instr_write_data[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput471 net471 instr_write_data[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput482 net482 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput493 net493 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output418_I net418 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_170_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0478__I3 _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_147_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0883__I0 net489 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1200_ net35 net464 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1093__CLK net681 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_239_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1062_ _0191_ _0153_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_230_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0874__I0 net421 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_202_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0915_ net488 net55 _0054_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0846_ net16 net149 _0436_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0777_ _0397_ net559 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input149_I la_data_in[70] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input316_I uP_data_mem_addr[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_246_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_224_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0865__I0 net417 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_142_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_146_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_107_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1034__A3 _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_240_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0700_ _0354_ net591 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_11526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0784__A2 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0631_ _0295_ net425 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_9260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0562_ _0256_ net454 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_8570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0493_ _0208_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_7880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1045_ _0138_ _0141_ _0142_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_241_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_224_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0829_ _0427_ net583 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input266_I la_oenb[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output485_I net485 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0518__A2 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_229_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0614_ net37 net335 _0284_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_10655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_fanout683_I net684 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout708 net709 net708 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0545_ _0246_ net422 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0476_ net40 _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_230_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1028_ net697 _0114_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input383_I wbs_dat_i[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input77_I la_data_in[120] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0684__A1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_224_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0987__A2 _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput360 wbs_adr_i[24] net360 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput371 wbs_adr_i[5] net371 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_5582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput382 wbs_dat_i[14] net382 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput393 wbs_dat_i[24] net393 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_203_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0528_ data_load_addr\[1\] _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_0459_ _0176_ _0180_ _0171_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input131_I la_data_in[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input229_I la_oenb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_104_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_235_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput190 la_oenb[108] net190 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_3_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input179_I la_data_in[98] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput620 net620 la_data_out[96] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput631 net631 uP_instr[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_173_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput642 net642 uP_instr[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput653 net653 wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_236_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput664 net664 wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput675 net675 wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_216_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input346_I wbs_adr_i[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1064__A1 _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1055__A1 data_load_addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0931_ _0182_ net62 _0064_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0862_ _0026_ net599 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_239_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0793_ _0406_ net566 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_244_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1046__A1 _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input296_I la_oenb[89] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput450 net450 instr_mem_addr[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput461 net461 instr_write_data[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput472 net472 instr_write_data[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_212_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput483 net483 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_236_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput494 net494 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1037__A1 _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1061_ _0242_ _0151_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_168_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1028__A1 net697 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0614__S _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0914_ _0056_ net623 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_239_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0845_ _0425_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_176_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0776_ net116 _0396_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_100_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_245_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input211_I la_oenb[127] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input309_I uP_data_mem_addr[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_222_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_240_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_8015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output430_I net430 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_11549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0630_ net697 net327 _0294_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_10815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0561_ instr_load_addr\[5\] net323 _0252_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_8560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0492_ _0207_ net52 _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_193_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0792__I0 net432 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0609__S _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1044_ _0173_ _0139_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0828_ net8 net140 _0426_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_198_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0759_ _0376_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_217_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input161_I la_data_in[81] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input259_I la_oenb[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input22_I instr[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0535__I0 data_load_addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0988__I _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0526__I0 _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0613_ _0285_ net432 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_236_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_0544_ data_load_addr\[6\] net315 _0245_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_8390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout709 net710 net709 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_214_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout676_I net677 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_171_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0475_ _0193_ net494 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1027_ instr_load_addr\[10\] _0127_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_207_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input376_I wbs_cyc_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0684__A2 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0712__S _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput350 wbs_adr_i[15] net350 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput361 wbs_adr_i[25] net361 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput372 wbs_adr_i[6] net372 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput383 wbs_dat_i[15] net383 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_40_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput394 wbs_dat_i[25] net394 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_770 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_4871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_205_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1092__RN net705 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_11198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0738__I0 net641 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0527_ _0234_ net416 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0458_ net9 net26 _0177_ _0178_ _0166_ _0179_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_246_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input124_I la_data_in[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_3_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0977__I0 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1083__RN net707 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_219_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0729__I0 net637 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_210_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1162__I net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0593__A1 net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1074__RN net702 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_177_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_233_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput180 la_data_in[99] net180 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput191 la_oenb[109] net191 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_188_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0959__I0 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput610 net610 la_data_out[87] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_86_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0584__A1 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_153_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput621 net621 la_data_out[97] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput632 net632 uP_instr[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_160_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput643 net643 wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput654 net654 wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput665 net665 wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_67_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input241_I la_oenb[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input339_I uP_write_data[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_210_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output460_I net460 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_238_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1055__A2 data_load_addr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0930_ _0065_ net505 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0861_ net416 net156 _0022_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_200_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0792_ net432 net123 _0404_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_237_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1046__A2 _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input191_I la_oenb[109] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input289_I la_oenb[82] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input52_I io_in[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput440 net691 dataw_en vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput451 net451 instr_mem_addr[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput462 net462 instr_write_data[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_154_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput473 net690 instrw_en vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_216_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput484 net484 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput495 net495 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_233_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_196_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0720__S _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1060_ _0149_ _0151_ _0152_ _0154_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_210_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1028__A2 _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0913_ net487 net180 _0054_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0844_ _0435_ net590 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0775_ _0344_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0630__S _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1189_ net363 analog_io[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input204_I la_oenb[120] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_205_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1019__A2 _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0540__S _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output423_I net423 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1170__I net374 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0560_ _0255_ net453 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_9284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0491_ net51 _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_8594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0544__I1 net315 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_212_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1043_ _0231_ _0235_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_4_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0625__S _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_241_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0827_ _0425_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_235_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0758_ _0386_ net550 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0689_ _0343_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input154_I la_data_in[75] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input321_I uP_instr_mem_addr[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__0535__I1 net312 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input15_I data_read_data[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0999__A1 instr_load_addr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0535__S _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_161_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output638_I net638 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_192_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1165__I net369 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0526__I1 net309 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_10635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0612_ net36 net334 _0284_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_9070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0543_ _0244_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_234_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0474_ _0191_ _0192_ _0189_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_7690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input7_I data_read_data[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1026_ _0096_ _0125_ _0127_ _0128_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_165_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input271_I la_oenb[66] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_200_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input369_I wbs_adr_i[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output490_I net490 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_213_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_200_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput340 uP_write_data[8] net340 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_6296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput351 wbs_adr_i[16] net351 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput362 wbs_adr_i[26] net362 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput373 wbs_adr_i[7] net373 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_20_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput384 wbs_dat_i[16] net384 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_79_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_760 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xinput395 wbs_dat_i[26] net395 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_771 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_4872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0526_ _0231_ net309 _0233_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0457_ net52 _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input117_I la_data_in[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_97_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_182_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_108_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1009_ _0096_ _0111_ _0113_ _0115_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_162_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input82_I la_data_in[125] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_182_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0977__I1 net342 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput170 la_data_in[8] net170 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_40_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput181 la_data_in[9] net181 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput192 la_oenb[10] net192 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_fanout701_I net702 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_203_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput600 net600 la_data_out[78] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_192_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput611 net611 la_data_out[88] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_66_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput622 net622 la_data_out[98] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput633 net633 uP_instr[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput644 net644 wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_236_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput655 net655 wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput666 net666 wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0509_ instr_load_addr\[12\] _0203_ _0205_ net4 _0208_ net21 _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_210_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input234_I la_oenb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input401_I wbs_dat_i[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_8913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output453_I net453 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_234_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1173__I net346 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_228_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0638__I0 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_163_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0860_ _0025_ net598 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0791_ _0405_ net565 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_239_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0810__I0 net425 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_174_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_168_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0989_ _0173_ _0099_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input184_I la_oenb[102] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_195_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0801__I0 net436 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput430 net430 data_write_data[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput441 net441 dataw_en_8bit[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput452 net452 instr_mem_addr[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input351_I wbs_adr_i[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput463 net463 instr_write_data[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput474 net474 instrw_en_8bit[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_173_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput485 net485 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_input45_I io_in[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput496 net496 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_5_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_223_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1168__I net372 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout690 net473 net690 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_232_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0448__S _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_246_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0859__I0 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0912_ _0055_ net622 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_204_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0843_ net15 net147 _0431_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_200_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0774_ _0395_ net557 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_192_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_fanout699_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1257_ net401 net668 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1188_ net362 analog_io[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_4_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_228_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_209_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input399_I wbs_dat_i[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0821__S _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_8006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output416_I net416 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_240_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_193_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0490_ _0205_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_8595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1042_ _0231_ _0138_ _0140_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0826_ _0424_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0757_ net449 net107 _0382_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__0440__I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0688_ _0346_ net547 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input147_I la_data_in[69] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input314_I uP_data_mem_addr[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0999__A2 instr_load_addr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1181__I net354 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_229_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0611_ _0244_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_10625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0542_ net694 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_8370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0473_ net12 net29 data_load_addr\[5\] instr_load_addr\[5\] _0183_ _0179_ _0192_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_7680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0636__S _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1025_ net698 _0109_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_228_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0809_ _0415_ net574 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_239_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input264_I la_oenb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0546__S _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_187_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output483_I net483 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1176__I net349 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput330 uP_write_data[13] net330 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_231_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput341 uP_write_data[9] net341 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_188_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput352 wbs_adr_i[17] net352 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput363 wbs_adr_i[27] net363 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput374 wbs_adr_i[8] net374 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_750 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_236_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput385 wbs_dat_i[17] net385 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_761 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_4862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput396 wbs_dat_i[27] net396 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xio_interface_772 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_166_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_242_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0525_ _0232_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0456_ instr_load_addr\[2\] _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0520__B1 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_149_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_180_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_56_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1008_ _0191_ _0114_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input381_I wbs_dat_i[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_194_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input75_I la_data_in[119] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_198_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1000__A1 _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1067__A1 _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_196_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput160 la_data_in[80] net160 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_20_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput171 la_data_in[90] net171 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput182 la_oenb[100] net182 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_94_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput193 la_oenb[110] net193 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_242_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput601 net601 la_data_out[79] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_236_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput612 net612 la_data_out[89] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput623 net623 la_data_out[99] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput634 net634 uP_instr[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_233_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput645 net645 wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_86_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput656 net656 wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput667 net667 wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0508_ _0217_ _0218_ _0220_ net484 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input227_I la_oenb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_223_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1049__A1 _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0734__S _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_243_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1055__A4 data_load_addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0790_ net431 net122 _0404_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_220_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0443__I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0988_ _0094_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input177_I la_data_in[96] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput420 net420 data_mem_addr[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_82_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput431 net431 data_write_data[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput442 net442 dataw_en_8bit[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_216_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput453 net453 instr_mem_addr[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput464 net464 instr_write_data[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput475 net475 instrw_en_8bit[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput486 net486 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_236_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input344_I wbs_adr_i[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput497 net497 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_87_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input38_I io_in[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0819__S _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1086__CLK net685 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1184__I net358 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout680 net684 net680 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_130_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout691 net693 net691 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_1_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0528__I data_load_addr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0464__S _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0911_ net486 net179 _0054_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_230_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0842_ _0434_ net589 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0773_ net456 net114 _0392_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_211_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1256_ net400 net667 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1187_ net361 analog_io[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_4_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input294_I la_oenb[87] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_220_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0901__I _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_218_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0786__I0 net424 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0549__S _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_216_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0710__I0 net367 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1179__I net352 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_8585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0529__I0 _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0459__S _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_232_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1041_ _0164_ _0139_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_219_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0701__I0 net414 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0825_ _0343_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0756_ _0385_ net549 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_213_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0687_ net104 _0345_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_157_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1239_ net381 net648 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input307_I la_oenb[99] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0687__A2 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0931__I0 _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0610_ _0283_ net431 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_10626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0541_ _0243_ net421 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_9094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_218_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0472_ net39 _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0922__I0 _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1024_ _0120_ _0126_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_223_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0808_ net439 net131 _0414_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_217_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0739_ _0375_ net541 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input257_I la_oenb[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input20_I instr[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0913__I0 net487 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_190_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output643_I net643 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1192__I net691 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput320 uP_instr_mem_addr[2] net320 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_6276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput331 uP_write_data[14] net331 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_213_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput342 wb_clk_i net342 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput353 wbs_adr_i[18] net353 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0904__I0 net483 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput364 wbs_adr_i[28] net364 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xio_interface_740 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_229_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput375 wbs_adr_i[9] net375 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_751 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput386 wbs_dat_i[18] net386 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_762 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xinput397 wbs_dat_i[28] net397 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_773 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_131_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0524_ net694 _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_8190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0455_ data_load_addr\[2\] _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0520__A1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0520__B2 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_208_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0446__I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_169_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1007_ _0093_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_219_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input374_I wbs_adr_i[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_191_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input68_I la_data_in[112] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1000__A2 _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_10990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1187__I net361 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput150 la_data_in[71] net150 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput161 la_data_in[81] net161 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput172 la_data_in[91] net172 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput183 la_oenb[101] net183 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput194 la_oenb[111] net194 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0569__A1 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_173_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput602 net602 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput613 net613 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput624 net624 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_10253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput635 net635 uP_instr[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput646 net646 wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput657 net657 wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput668 net668 wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0507_ _0219_ net696 _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_228_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input122_I la_data_in[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output439_I net439 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_172_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0987_ _0248_ _0250_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_220_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput421 net421 data_mem_addr[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_172_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput432 net432 data_write_data[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput443 net443 dataw_en_8bit[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput454 net454 instr_mem_addr[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput465 net465 instr_write_data[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput476 net476 instrw_en_8bit[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput487 net487 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput498 net498 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_160_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input337_I uP_write_data[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout681 net683 net681 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_219_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout692 net693 net692 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_21_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0910_ _0048_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_0841_ net14 net146 _0431_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_239_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0772_ _0394_ net556 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_237_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1255_ net398 net665 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1186_ net360 analog_io[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_25_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_224_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0454__I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0483__I0 _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_222_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input287_I la_oenb[80] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_229_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input50_I io_in[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0474__I0 _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_240_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_11509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_9232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1195__I net692 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0529__I1 net310 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_7885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1040_ _0137_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0824_ _0423_ net582 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0755_ net633 net106 _0382_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_200_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0686_ _0344_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_171_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1238_ net380 net647 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1169_ net373 analog_io[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input202_I la_oenb[119] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0999__A4 instr_load_addr\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_146_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input98_I la_data_in[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_165_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output421_I net421 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0695__I0 net411 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_200_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0540_ _0242_ net314 _0238_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_9095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_8361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0471_ _0190_ net493 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_7660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1023_ instr_load_addr\[8\] instr_load_addr\[9\] _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_241_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__0933__S _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_245_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0807_ _0403_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_219_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0738_ net641 net98 _0371_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_232_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0669_ net264 net253 net286 net275 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_193_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input152_I la_data_in[73] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input13_I data_read_data[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_233_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output469_I net469 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output636_I net636 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_6211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput310 uP_data_mem_addr[1] net310 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_153_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput321 uP_instr_mem_addr[3] net321 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_6277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput332 uP_write_data[15] net332 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_6288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput343 wb_rst_i net343 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput354 wbs_adr_i[19] net354 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_730 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput365 wbs_adr_i[29] net365 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xio_interface_741 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_188_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput376 wbs_cyc_i net376 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_752 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_40_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput387 wbs_dat_i[19] net387 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_763 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_5_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput398 wbs_dat_i[29] net398 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_774 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_4875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_203_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0523_ data_load_addr\[0\] _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_8180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0454_ net36 _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_7490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I data_read_data[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__0520__A2 _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_215_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1006_ _0107_ _0112_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_126_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_9809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input367_I wbs_adr_i[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_210_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__0898__I0 net497 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput140 la_data_in[62] net140 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_42_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput151 la_data_in[72] net151 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_98_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput162 la_data_in[82] net162 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0889__I0 net493 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput173 la_data_in[92] net173 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput184 la_oenb[102] net184 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput195 la_oenb[112] net195 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__0502__A2 net697 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0483__S _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_220_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput603 net603 la_data_out[80] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_86_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput614 net614 la_data_out[90] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_236_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput625 net625 reset vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput636 net636 uP_instr[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput647 net647 wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput658 net658 wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput669 net669 wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_64_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_116_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0506_ _0201_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0457__I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_228_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input115_I la_data_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input80_I la_data_in[123] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_9617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_191_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1198__I net440 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_209_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0986_ _0248_ _0095_ _0097_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0740__I _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_145_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput422 net422 data_mem_addr[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput433 net433 data_write_data[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput444 net444 dataw_en_8bit[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput455 net455 instr_mem_addr[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput466 net466 instr_write_data[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput477 net477 instrw_en_8bit[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_216_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput488 net488 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_233_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput499 net499 la_data_out[100] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_232_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0714__A2 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input232_I la_oenb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output451_I net451 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_8757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout682 net683 net682 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout693 net440 net693 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_4_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0840_ _0433_ net588 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0771_ net455 net113 _0392_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1254_ net397 net664 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1185_ net359 analog_io[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_98_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_221_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0969_ net317 net80 _0085_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input182_I la_oenb[100] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input43_I io_in[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_5906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_9277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_9299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0823_ net1 net139 _0419_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0754_ _0384_ net548 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__0473__S0 _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout697_I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_0685_ _0343_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1237_ net379 net646 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1168_ net372 analog_io[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input397_I wbs_dat_i[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1030__A1 instr_load_addr\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_194_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_7138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_7149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_240_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_221_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_9052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_9085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_9096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_8351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_8362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_8384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_0470_ _0186_ _0188_ _0189_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_234_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_7650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_7661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_7694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1022_ instr_load_addr\[8\] _0121_ instr_load_addr\[9\] _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_241_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0806_ _0413_ net573 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1012__A1 _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0737_ _0374_ net540 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_217_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0668_ net242 net231 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_0599_ net22 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input145_I la_data_in[67] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_4309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input312_I uP_data_mem_addr[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_226_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_228_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1020__S _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_224_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output629_I net629 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_235_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput300 la_oenb[92] net300 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput311 uP_data_mem_addr[2] net311 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_216_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput322 uP_instr_mem_addr[4] net322 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_131_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput333 uP_write_data[1] net333 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_6289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput344 wbs_adr_i[0] net344 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_720 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__0514__B1 _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_188_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput355 wbs_adr_i[1] net355 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xio_interface_731 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput366 wbs_adr_i[2] net366 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_4832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_742 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_131_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput377 wbs_dat_i[0] net377 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput388 wbs_dat_i[1] net388 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xio_interface_753 irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_79_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_764 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xinput399 wbs_dat_i[2] net399 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xio_interface_775 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_4876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_11104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_200_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_11115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_11137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_11159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_0522_ _0211_ _0229_ _0230_ net488 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_153_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_8181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_8192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0453_ _0175_ net489 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_7480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_7491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__0505__C2 net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1005_ instr_load_addr\[4\] instr_load_addr\[5\] _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_225_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input262_I la_oenb[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_10970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1089__CLK net677 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output481_I net481 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_210_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput130 la_data_in[53] net130 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput141 la_data_in[63] net141 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_24_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput152 la_data_in[73] net152 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput163 la_data_in[83] net163 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput174 la_data_in[93] net174 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput185 la_oenb[103] net185 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_94_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput196 la_oenb[113] net196 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_4662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_10211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_10222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput604 net604 la_data_out[81] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput615 net615 la_data_out[91] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_10244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_10255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput626 net626 start vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput637 net637 uP_instr[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_233_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput648 net648 wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_99_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput659 net659 wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_47_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_10288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_10299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_0505_ instr_load_addr\[11\] _0204_ _0206_ net3 _0209_ net20 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_236_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
.ends

