// This is the unpowered netlist.
module matrix_multiply (clk,
    execute,
    reset,
    input_val,
    result,
    sel_in,
    sel_out);
 input clk;
 input execute;
 input reset;
 input [7:0] input_val;
 output [16:0] result;
 input [2:0] sel_in;
 input [1:0] sel_out;

 wire \A[0][0] ;
 wire \A[0][1] ;
 wire \A[0][2] ;
 wire \A[0][3] ;
 wire \A[0][4] ;
 wire \A[0][5] ;
 wire \A[0][6] ;
 wire \A[0][7] ;
 wire \A[1][0] ;
 wire \A[1][1] ;
 wire \A[1][2] ;
 wire \A[1][3] ;
 wire \A[1][4] ;
 wire \A[1][5] ;
 wire \A[1][6] ;
 wire \A[1][7] ;
 wire \A[2][0] ;
 wire \A[2][1] ;
 wire \A[2][2] ;
 wire \A[2][3] ;
 wire \A[2][4] ;
 wire \A[2][5] ;
 wire \A[2][6] ;
 wire \A[2][7] ;
 wire \A[3][0] ;
 wire \A[3][1] ;
 wire \A[3][2] ;
 wire \A[3][3] ;
 wire \A[3][4] ;
 wire \A[3][5] ;
 wire \A[3][6] ;
 wire \A[3][7] ;
 wire \B[0][0] ;
 wire \B[0][1] ;
 wire \B[0][2] ;
 wire \B[0][3] ;
 wire \B[0][4] ;
 wire \B[0][5] ;
 wire \B[0][6] ;
 wire \B[0][7] ;
 wire \B[1][0] ;
 wire \B[1][1] ;
 wire \B[1][2] ;
 wire \B[1][3] ;
 wire \B[1][4] ;
 wire \B[1][5] ;
 wire \B[1][6] ;
 wire \B[1][7] ;
 wire \B[2][0] ;
 wire \B[2][1] ;
 wire \B[2][2] ;
 wire \B[2][3] ;
 wire \B[2][4] ;
 wire \B[2][5] ;
 wire \B[2][6] ;
 wire \B[2][7] ;
 wire \B[3][0] ;
 wire \B[3][1] ;
 wire \B[3][2] ;
 wire \B[3][3] ;
 wire \B[3][4] ;
 wire \B[3][5] ;
 wire \B[3][6] ;
 wire \B[3][7] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;

 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3400_ (.I(net15),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3401_ (.A1(net16),
    .A2(_0674_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3402_ (.I(_0685_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3403_ (.I(\B[3][6] ),
    .Z(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3404_ (.I(\A[3][0] ),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3405_ (.A1(_0707_),
    .A2(_0718_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3406_ (.I(\A[3][2] ),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3407_ (.I(\B[3][4] ),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3408_ (.A1(_0740_),
    .A2(_0751_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3409_ (.I(\B[3][5] ),
    .Z(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3410_ (.A1(_0773_),
    .A2(\A[3][1] ),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3411_ (.A1(_0762_),
    .A2(_0784_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3412_ (.A1(_0729_),
    .A2(_0795_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3413_ (.I(\B[3][2] ),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3414_ (.I(\A[3][4] ),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3415_ (.A1(_0817_),
    .A2(_0828_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3416_ (.I(\B[3][1] ),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3417_ (.I(_0850_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3418_ (.I(\A[3][3] ),
    .Z(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3419_ (.I(_0872_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3420_ (.A1(_0861_),
    .A2(_0883_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3421_ (.I(_0740_),
    .Z(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3422_ (.I(\B[3][3] ),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3423_ (.I(_0916_),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3424_ (.A1(_0905_),
    .A2(_0927_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3425_ (.I(\B[3][2] ),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3426_ (.I(_0949_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3427_ (.I(_0960_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3428_ (.I(_0872_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3429_ (.I(_0828_),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3430_ (.I(_0850_),
    .Z(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3431_ (.I(_1004_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3432_ (.A1(_0971_),
    .A2(_0982_),
    .B1(_0993_),
    .B2(_1015_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3433_ (.A1(_0839_),
    .A2(_0894_),
    .B1(_0938_),
    .B2(_1026_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3434_ (.I(\A[3][5] ),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3435_ (.A1(_1048_),
    .A2(_0850_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3436_ (.I(\A[3][3] ),
    .Z(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3437_ (.I(\B[3][3] ),
    .Z(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3438_ (.A1(_1070_),
    .A2(_1081_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3439_ (.A1(_1059_),
    .A2(_0839_),
    .A3(_1092_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3440_ (.A1(_1037_),
    .A2(_1103_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3441_ (.A1(_1037_),
    .A2(_1103_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3442_ (.A1(_0806_),
    .A2(_1114_),
    .B(_1125_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3443_ (.I(\A[2][2] ),
    .Z(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3444_ (.I(\B[1][3] ),
    .Z(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3445_ (.A1(_1147_),
    .A2(_1158_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3446_ (.I(\A[2][1] ),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3447_ (.I(\B[1][4] ),
    .Z(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3448_ (.A1(_1180_),
    .A2(_1191_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3449_ (.A1(_1169_),
    .A2(_1202_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3450_ (.I(\B[1][5] ),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3451_ (.I(_1224_),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3452_ (.I(\A[2][0] ),
    .Z(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3453_ (.A1(_1235_),
    .A2(_1246_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3454_ (.A1(_1169_),
    .A2(_1202_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3455_ (.A1(_1257_),
    .A2(_1268_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3456_ (.I(\B[1][6] ),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3457_ (.I(_1290_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3458_ (.I(_1301_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3459_ (.I(_1246_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3460_ (.A1(_1312_),
    .A2(_1323_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3461_ (.I(\A[3][6] ),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3462_ (.I(_1345_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3463_ (.I(_1356_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3464_ (.I(_1367_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3465_ (.I(\B[3][0] ),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3466_ (.A1(_1378_),
    .A2(_1389_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3467_ (.A1(_1334_),
    .A2(_1400_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3468_ (.A1(_1334_),
    .A2(_1400_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3469_ (.A1(_1213_),
    .A2(_1279_),
    .B(_1411_),
    .C(_1422_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3470_ (.I(\A[3][5] ),
    .Z(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3471_ (.A1(_1444_),
    .A2(_0817_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3472_ (.A1(_0861_),
    .A2(_0993_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3473_ (.A1(_1059_),
    .A2(_0839_),
    .Z(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3474_ (.A1(_1455_),
    .A2(_1466_),
    .B1(_1092_),
    .B2(_1477_),
    .ZN(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3475_ (.I(\A[3][6] ),
    .Z(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3476_ (.I(\B[3][1] ),
    .Z(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3477_ (.A1(_1499_),
    .A2(_1510_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3478_ (.I(\A[3][4] ),
    .Z(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3479_ (.A1(_1081_),
    .A2(_1532_),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3480_ (.A1(_1521_),
    .A2(_1455_),
    .A3(_1543_),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3481_ (.I(\B[3][6] ),
    .Z(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3482_ (.I(\A[3][1] ),
    .Z(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3483_ (.A1(_1565_),
    .A2(_1576_),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3484_ (.I(\B[3][4] ),
    .Z(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3485_ (.A1(_0872_),
    .A2(_1598_),
    .ZN(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3486_ (.I(\B[3][5] ),
    .Z(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3487_ (.A1(_1620_),
    .A2(_0740_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3488_ (.A1(_1609_),
    .A2(_1631_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3489_ (.A1(_1587_),
    .A2(_1642_),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3490_ (.A1(_1488_),
    .A2(_1554_),
    .A3(_1653_),
    .Z(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3491_ (.A1(_1433_),
    .A2(_1664_),
    .Z(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3492_ (.A1(_1433_),
    .A2(_1664_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3493_ (.A1(_1136_),
    .A2(_1675_),
    .B(_1686_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3494_ (.A1(_1620_),
    .A2(_0872_),
    .ZN(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3495_ (.A1(_1708_),
    .A2(_0762_),
    .ZN(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3496_ (.A1(_1587_),
    .A2(_1642_),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3497_ (.A1(_1719_),
    .A2(_1730_),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3498_ (.A1(_1697_),
    .A2(_1741_),
    .Z(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3499_ (.A1(_1697_),
    .A2(_1741_),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3500_ (.A1(_1752_),
    .A2(_1763_),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3501_ (.I(\B[3][7] ),
    .Z(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3502_ (.I(_1576_),
    .Z(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3503_ (.I(_1796_),
    .Z(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3504_ (.I(_1807_),
    .Z(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3505_ (.I(_1818_),
    .Z(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3506_ (.A1(_1785_),
    .A2(_1829_),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3507_ (.A1(_1774_),
    .A2(_1840_),
    .Z(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3508_ (.A1(_1136_),
    .A2(_1675_),
    .Z(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3509_ (.I(_1862_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3510_ (.A1(_1213_),
    .A2(_1279_),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3511_ (.A1(_1422_),
    .A2(_1411_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3512_ (.A1(_1883_),
    .A2(_1894_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3513_ (.A1(_1257_),
    .A2(_1268_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3514_ (.I(\B[1][1] ),
    .Z(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3515_ (.I(_1927_),
    .Z(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3516_ (.I(\A[2][4] ),
    .Z(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3517_ (.A1(_1938_),
    .A2(_1949_),
    .ZN(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3518_ (.I(\B[1][0] ),
    .Z(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3519_ (.I(_1971_),
    .Z(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3520_ (.I(\A[2][3] ),
    .Z(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3521_ (.I(_1993_),
    .Z(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3522_ (.A1(_1982_),
    .A2(_2004_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3523_ (.I(_1147_),
    .Z(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3524_ (.I(\B[1][2] ),
    .Z(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3525_ (.I(_2037_),
    .Z(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3526_ (.A1(_2026_),
    .A2(_2048_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3527_ (.I(_1938_),
    .Z(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3528_ (.I(\A[2][4] ),
    .Z(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3529_ (.I(_2081_),
    .Z(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3530_ (.I(\B[1][0] ),
    .Z(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3531_ (.I(_2102_),
    .Z(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3532_ (.A1(_2070_),
    .A2(_2004_),
    .B1(_2092_),
    .B2(_2113_),
    .ZN(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3533_ (.A1(_1960_),
    .A2(_2015_),
    .B1(_2059_),
    .B2(_2124_),
    .ZN(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3534_ (.I(\A[2][5] ),
    .Z(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3535_ (.I(_2146_),
    .Z(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3536_ (.I(\B[1][0] ),
    .Z(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3537_ (.A1(_2157_),
    .A2(_2168_),
    .ZN(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3538_ (.I(\A[2][3] ),
    .Z(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3539_ (.I(_2190_),
    .Z(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3540_ (.A1(_2048_),
    .A2(_2201_),
    .ZN(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3541_ (.A1(_2179_),
    .A2(_1960_),
    .A3(_2212_),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3542_ (.A1(_2135_),
    .A2(_2223_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3543_ (.A1(_2135_),
    .A2(_2223_),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3544_ (.A1(_1916_),
    .A2(_2234_),
    .B(_2245_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3545_ (.I(_2190_),
    .Z(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3546_ (.A1(_2267_),
    .A2(_1158_),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3547_ (.I(\A[2][2] ),
    .Z(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3548_ (.I(\B[1][4] ),
    .Z(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3549_ (.I(_2299_),
    .Z(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3550_ (.A1(_2288_),
    .A2(_2310_),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3551_ (.I(\B[1][5] ),
    .Z(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3552_ (.I(_2332_),
    .Z(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3553_ (.I(\A[2][1] ),
    .Z(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3554_ (.A1(_2343_),
    .A2(_2354_),
    .ZN(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3555_ (.A1(_2277_),
    .A2(_2321_),
    .A3(_2365_),
    .Z(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3556_ (.I(\A[2][5] ),
    .Z(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3557_ (.I(\B[1][1] ),
    .Z(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3558_ (.A1(_2387_),
    .A2(_2398_),
    .ZN(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3559_ (.I(_2102_),
    .Z(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3560_ (.I(_2081_),
    .Z(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3561_ (.A1(_2419_),
    .A2(_2430_),
    .ZN(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3562_ (.I(_2387_),
    .Z(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3563_ (.A1(_2452_),
    .A2(_2419_),
    .B1(_2070_),
    .B2(_2430_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3564_ (.A1(_2408_),
    .A2(_2441_),
    .B1(_2212_),
    .B2(_2463_),
    .ZN(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3565_ (.I(\B[1][2] ),
    .Z(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3566_ (.I(\A[2][4] ),
    .Z(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3567_ (.A1(_2484_),
    .A2(_2495_),
    .ZN(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3568_ (.I(\A[2][6] ),
    .Z(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3569_ (.I(_2515_),
    .Z(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3570_ (.A1(_2525_),
    .A2(_1971_),
    .ZN(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3571_ (.A1(_2408_),
    .A2(_2505_),
    .A3(_2535_),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3572_ (.A1(_2473_),
    .A2(_2545_),
    .ZN(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3573_ (.A1(_2376_),
    .A2(_2555_),
    .Z(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3574_ (.A1(_2256_),
    .A2(_2565_),
    .Z(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3575_ (.A1(_2256_),
    .A2(_2565_),
    .Z(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3576_ (.A1(_1905_),
    .A2(_2576_),
    .B(_2586_),
    .ZN(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3577_ (.A1(_2473_),
    .A2(_2545_),
    .ZN(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3578_ (.A1(_2376_),
    .A2(_2555_),
    .B(_2606_),
    .ZN(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3579_ (.A1(_1993_),
    .A2(_1191_),
    .ZN(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3580_ (.A1(_1224_),
    .A2(_1147_),
    .ZN(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3581_ (.I(\B[1][3] ),
    .Z(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3582_ (.I(_2644_),
    .Z(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3583_ (.I(_1949_),
    .Z(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3584_ (.A1(_2651_),
    .A2(_2660_),
    .ZN(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3585_ (.A1(_2627_),
    .A2(_2636_),
    .A3(_2668_),
    .Z(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3586_ (.A1(\A[2][6] ),
    .A2(_1927_),
    .ZN(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3587_ (.I(\A[2][6] ),
    .Z(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3588_ (.I(_1927_),
    .Z(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3589_ (.I(_2146_),
    .Z(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3590_ (.A1(_2690_),
    .A2(_2102_),
    .B1(_2697_),
    .B2(_2704_),
    .ZN(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3591_ (.A1(_2179_),
    .A2(_2684_),
    .B1(_2711_),
    .B2(_2505_),
    .ZN(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3592_ (.A1(_2146_),
    .A2(_2484_),
    .ZN(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3593_ (.I(\A[2][7] ),
    .Z(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3594_ (.A1(_2732_),
    .A2(_2168_),
    .ZN(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3595_ (.A1(_2684_),
    .A2(_2725_),
    .A3(_2739_),
    .ZN(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3596_ (.A1(_2718_),
    .A2(_2746_),
    .ZN(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3597_ (.A1(_2676_),
    .A2(_2753_),
    .Z(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3598_ (.A1(_2277_),
    .A2(_2321_),
    .Z(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3599_ (.A1(_2627_),
    .A2(_1169_),
    .B1(_2365_),
    .B2(_2758_),
    .ZN(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3600_ (.I(\A[3][7] ),
    .Z(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3601_ (.A1(_2760_),
    .A2(_1389_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3602_ (.I(\B[1][6] ),
    .Z(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3603_ (.I(\B[1][7] ),
    .Z(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3604_ (.A1(_2762_),
    .A2(_2763_),
    .A3(\A[2][0] ),
    .A4(\A[2][1] ),
    .Z(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3605_ (.I(\B[1][7] ),
    .Z(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3606_ (.I(_2765_),
    .Z(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3607_ (.A1(_2766_),
    .A2(\A[2][0] ),
    .B1(_1180_),
    .B2(_1290_),
    .ZN(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3608_ (.A1(_2761_),
    .A2(_2764_),
    .A3(_2767_),
    .Z(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3609_ (.A1(_2764_),
    .A2(_2767_),
    .B(_2761_),
    .ZN(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3610_ (.A1(_2768_),
    .A2(_2769_),
    .Z(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3611_ (.A1(_2759_),
    .A2(_2770_),
    .ZN(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3612_ (.A1(_1422_),
    .A2(_2771_),
    .ZN(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3613_ (.A1(_2616_),
    .A2(_2757_),
    .A3(_2772_),
    .ZN(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3614_ (.A1(_2596_),
    .A2(_2773_),
    .Z(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3615_ (.A1(_1905_),
    .A2(_2576_),
    .Z(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3616_ (.A1(_2586_),
    .A2(_2775_),
    .B(_2773_),
    .ZN(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3617_ (.A1(_1872_),
    .A2(_2774_),
    .B(_2776_),
    .ZN(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3618_ (.A1(_2759_),
    .A2(_2770_),
    .ZN(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3619_ (.A1(_1422_),
    .A2(_2771_),
    .B(_2778_),
    .ZN(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3620_ (.A1(_0707_),
    .A2(_0905_),
    .ZN(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3621_ (.A1(_1532_),
    .A2(_1598_),
    .ZN(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3622_ (.A1(_2781_),
    .A2(_1708_),
    .ZN(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3623_ (.A1(_2780_),
    .A2(_2782_),
    .ZN(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3624_ (.A1(_1345_),
    .A2(_0949_),
    .ZN(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3625_ (.I(_1499_),
    .Z(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3626_ (.I(_0817_),
    .Z(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3627_ (.I(_1444_),
    .Z(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3628_ (.A1(_2785_),
    .A2(_0861_),
    .B1(_2786_),
    .B2(_2787_),
    .ZN(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3629_ (.A1(_2784_),
    .A2(_1059_),
    .B1(_1543_),
    .B2(_2788_),
    .ZN(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3630_ (.I(\A[3][7] ),
    .Z(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3631_ (.A1(_2790_),
    .A2(_0850_),
    .ZN(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3632_ (.A1(_1048_),
    .A2(_0916_),
    .ZN(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3633_ (.A1(_2784_),
    .A2(_2791_),
    .A3(_2792_),
    .ZN(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3634_ (.A1(_2789_),
    .A2(_2793_),
    .ZN(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3635_ (.A1(_2783_),
    .A2(_2794_),
    .Z(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3636_ (.A1(_1488_),
    .A2(_1554_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3637_ (.A1(_1488_),
    .A2(_1554_),
    .ZN(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3638_ (.A1(_1653_),
    .A2(_2796_),
    .B(_2797_),
    .ZN(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3639_ (.A1(_2779_),
    .A2(_2795_),
    .A3(_2798_),
    .ZN(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3640_ (.A1(_2616_),
    .A2(_2757_),
    .ZN(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3641_ (.A1(_2616_),
    .A2(_2757_),
    .ZN(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3642_ (.A1(_2772_),
    .A2(_2800_),
    .B(_2801_),
    .ZN(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3643_ (.A1(_2761_),
    .A2(_2764_),
    .A3(_2767_),
    .ZN(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3644_ (.A1(_2764_),
    .A2(_2803_),
    .ZN(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3645_ (.A1(_2495_),
    .A2(_2299_),
    .ZN(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3646_ (.I(_2190_),
    .Z(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3647_ (.A1(_2651_),
    .A2(_2660_),
    .B1(_2310_),
    .B2(_2806_),
    .ZN(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3648_ (.A1(_2277_),
    .A2(_2805_),
    .B1(_2807_),
    .B2(_2636_),
    .ZN(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3649_ (.I(_2763_),
    .Z(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3650_ (.I(_1147_),
    .Z(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3651_ (.A1(_2809_),
    .A2(_2354_),
    .B1(_2810_),
    .B2(_1301_),
    .ZN(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3652_ (.I(_2762_),
    .Z(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3653_ (.I(_2765_),
    .Z(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3654_ (.I(\A[2][1] ),
    .Z(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3655_ (.A1(_2812_),
    .A2(_2813_),
    .A3(_2814_),
    .A4(_2288_),
    .Z(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3656_ (.A1(_2811_),
    .A2(_2815_),
    .ZN(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3657_ (.A1(_2808_),
    .A2(_2816_),
    .Z(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3658_ (.A1(_2804_),
    .A2(_2817_),
    .Z(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3659_ (.A1(_2718_),
    .A2(_2746_),
    .ZN(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3660_ (.A1(_2676_),
    .A2(_2753_),
    .B(_2819_),
    .ZN(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3661_ (.I(\A[2][6] ),
    .Z(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3662_ (.A1(_2732_),
    .A2(_2168_),
    .B1(_1938_),
    .B2(_2821_),
    .ZN(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3663_ (.A1(_2732_),
    .A2(_2821_),
    .A3(_2168_),
    .A4(_2398_),
    .ZN(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3664_ (.A1(_2725_),
    .A2(_2822_),
    .B(_2823_),
    .ZN(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3665_ (.A1(\A[2][7] ),
    .A2(_1927_),
    .ZN(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3666_ (.A1(_2515_),
    .A2(_2484_),
    .ZN(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3667_ (.A1(_2825_),
    .A2(_2826_),
    .Z(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3668_ (.A1(_2824_),
    .A2(_2827_),
    .ZN(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3669_ (.A1(_2387_),
    .A2(\B[1][3] ),
    .ZN(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3670_ (.A1(_1224_),
    .A2(_1993_),
    .ZN(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3671_ (.A1(_2805_),
    .A2(_2829_),
    .A3(_2830_),
    .Z(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3672_ (.A1(_2828_),
    .A2(_2831_),
    .Z(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3673_ (.A1(_2820_),
    .A2(_2832_),
    .ZN(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3674_ (.A1(_2818_),
    .A2(_2833_),
    .Z(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3675_ (.A1(_2802_),
    .A2(_2834_),
    .ZN(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3676_ (.A1(_2799_),
    .A2(_2835_),
    .Z(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3677_ (.A1(_2777_),
    .A2(_2836_),
    .Z(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3678_ (.A1(_2777_),
    .A2(_2836_),
    .Z(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3679_ (.A1(_1851_),
    .A2(_2837_),
    .B(_2838_),
    .ZN(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3680_ (.A1(_2779_),
    .A2(_2795_),
    .Z(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3681_ (.A1(_2779_),
    .A2(_2795_),
    .Z(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3682_ (.A1(_2798_),
    .A2(_2840_),
    .B(_2841_),
    .ZN(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3683_ (.A1(\B[3][5] ),
    .A2(\A[3][4] ),
    .ZN(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3684_ (.A1(_1609_),
    .A2(_2843_),
    .ZN(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3685_ (.A1(_2780_),
    .A2(_2782_),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3686_ (.A1(_2844_),
    .A2(_2845_),
    .ZN(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3687_ (.A1(_2842_),
    .A2(_2846_),
    .Z(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3688_ (.I(_0905_),
    .Z(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3689_ (.I(_2848_),
    .Z(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3690_ (.A1(_1785_),
    .A2(_2849_),
    .ZN(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3691_ (.A1(_2847_),
    .A2(_2850_),
    .ZN(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3692_ (.A1(_2802_),
    .A2(_2834_),
    .ZN(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3693_ (.A1(_2799_),
    .A2(_2835_),
    .B(_2852_),
    .ZN(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3694_ (.A1(_2783_),
    .A2(_2794_),
    .ZN(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3695_ (.A1(_2789_),
    .A2(_2793_),
    .B(_2854_),
    .ZN(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3696_ (.A1(_2808_),
    .A2(_2816_),
    .ZN(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3697_ (.A1(_2808_),
    .A2(_2816_),
    .ZN(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3698_ (.A1(_2804_),
    .A2(_2856_),
    .B(_2857_),
    .ZN(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3699_ (.A1(_1565_),
    .A2(_1070_),
    .ZN(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3700_ (.A1(_1444_),
    .A2(\B[3][4] ),
    .ZN(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3701_ (.A1(_2843_),
    .A2(_2860_),
    .ZN(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3702_ (.A1(_2859_),
    .A2(_2861_),
    .ZN(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3703_ (.I(_0949_),
    .Z(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3704_ (.A1(_2760_),
    .A2(_1510_),
    .B1(_2863_),
    .B2(_1499_),
    .ZN(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3705_ (.A1(_2760_),
    .A2(_1356_),
    .A3(_1510_),
    .A4(_2863_),
    .ZN(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3706_ (.A1(_2864_),
    .A2(_2792_),
    .B(_2865_),
    .ZN(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3707_ (.A1(\A[3][7] ),
    .A2(_0949_),
    .ZN(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3708_ (.A1(_1345_),
    .A2(_0916_),
    .ZN(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3709_ (.A1(_2867_),
    .A2(_2868_),
    .Z(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3710_ (.A1(_2866_),
    .A2(_2869_),
    .ZN(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3711_ (.A1(_2862_),
    .A2(_2870_),
    .Z(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3712_ (.A1(_2858_),
    .A2(_2871_),
    .ZN(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3713_ (.A1(_2855_),
    .A2(_2872_),
    .ZN(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3714_ (.A1(_2820_),
    .A2(_2832_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3715_ (.A1(_2818_),
    .A2(_2833_),
    .B(_2874_),
    .ZN(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3716_ (.A1(_2387_),
    .A2(\B[1][4] ),
    .ZN(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3717_ (.A1(_2805_),
    .A2(_2829_),
    .Z(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3718_ (.A1(_2668_),
    .A2(_2876_),
    .B1(_2877_),
    .B2(_2830_),
    .ZN(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3719_ (.I(_2765_),
    .Z(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3720_ (.A1(_2879_),
    .A2(_2288_),
    .ZN(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3721_ (.A1(_2812_),
    .A2(_2806_),
    .ZN(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3722_ (.I(\A[2][2] ),
    .Z(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3723_ (.A1(_1290_),
    .A2(_2766_),
    .A3(_2882_),
    .A4(_1993_),
    .Z(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3724_ (.A1(_2880_),
    .A2(_2881_),
    .B(_2883_),
    .ZN(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3725_ (.A1(_2878_),
    .A2(_2884_),
    .ZN(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3726_ (.A1(_2815_),
    .A2(_2885_),
    .Z(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3727_ (.A1(_2824_),
    .A2(_2827_),
    .ZN(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3728_ (.A1(_2828_),
    .A2(_2831_),
    .B(_2887_),
    .ZN(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3729_ (.A1(_2332_),
    .A2(_2495_),
    .ZN(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3730_ (.A1(_2690_),
    .A2(_2644_),
    .ZN(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3731_ (.A1(_2876_),
    .A2(_2889_),
    .A3(_2890_),
    .Z(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3732_ (.I(\A[2][7] ),
    .Z(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3733_ (.I(_2892_),
    .Z(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3734_ (.I(_2037_),
    .Z(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3735_ (.A1(_2893_),
    .A2(_2894_),
    .A3(_2684_),
    .ZN(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3736_ (.A1(_2891_),
    .A2(_2895_),
    .Z(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3737_ (.A1(_2888_),
    .A2(_2896_),
    .ZN(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3738_ (.A1(_2886_),
    .A2(_2897_),
    .Z(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3739_ (.A1(_2875_),
    .A2(_2898_),
    .ZN(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3740_ (.A1(_2873_),
    .A2(_2899_),
    .Z(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3741_ (.A1(_2853_),
    .A2(_2900_),
    .Z(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3742_ (.A1(_2851_),
    .A2(_2901_),
    .ZN(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3743_ (.A1(_2839_),
    .A2(_2902_),
    .ZN(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3744_ (.A1(_1774_),
    .A2(_1840_),
    .B(_1752_),
    .ZN(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3745_ (.A1(_2839_),
    .A2(_2902_),
    .Z(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3746_ (.A1(_2904_),
    .A2(_2905_),
    .Z(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3747_ (.I(\B[3][7] ),
    .Z(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3748_ (.I(_2907_),
    .Z(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3749_ (.I(_2908_),
    .Z(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3750_ (.I(_2849_),
    .Z(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3751_ (.A1(_2909_),
    .A2(_2910_),
    .A3(_2847_),
    .ZN(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3752_ (.A1(_2842_),
    .A2(_2846_),
    .B(_2911_),
    .ZN(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3753_ (.A1(_2853_),
    .A2(_2900_),
    .Z(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3754_ (.A1(_2851_),
    .A2(_2901_),
    .B(_2913_),
    .ZN(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3755_ (.A1(_2855_),
    .A2(_2872_),
    .ZN(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3756_ (.A1(_2858_),
    .A2(_2871_),
    .B(_2915_),
    .ZN(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3757_ (.A1(_2843_),
    .A2(_2860_),
    .ZN(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3758_ (.A1(_2859_),
    .A2(_2861_),
    .ZN(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3759_ (.A1(_2917_),
    .A2(_2918_),
    .ZN(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3760_ (.A1(_2916_),
    .A2(_2919_),
    .Z(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3761_ (.I(\B[3][7] ),
    .Z(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3762_ (.I(_0883_),
    .Z(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3763_ (.I(_2922_),
    .Z(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3764_ (.A1(_2921_),
    .A2(_2923_),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3765_ (.A1(_2920_),
    .A2(_2924_),
    .ZN(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3766_ (.A1(_2875_),
    .A2(_2898_),
    .ZN(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3767_ (.A1(_2873_),
    .A2(_2899_),
    .B(_2926_),
    .ZN(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3768_ (.A1(_2866_),
    .A2(_2869_),
    .ZN(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3769_ (.A1(_2862_),
    .A2(_2870_),
    .B(_2928_),
    .ZN(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3770_ (.I(_1312_),
    .Z(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3771_ (.I(_2814_),
    .Z(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3772_ (.I(_2931_),
    .Z(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3773_ (.I(_2932_),
    .Z(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3774_ (.A1(_2930_),
    .A2(_2933_),
    .ZN(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3775_ (.A1(_2878_),
    .A2(_2884_),
    .ZN(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3776_ (.A1(_2934_),
    .A2(_2880_),
    .A3(_2885_),
    .B(_2935_),
    .ZN(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3777_ (.I(_2790_),
    .Z(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3778_ (.I(_2937_),
    .Z(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3779_ (.I(_1081_),
    .Z(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3780_ (.I(_2939_),
    .Z(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3781_ (.A1(_2938_),
    .A2(_2940_),
    .A3(_2784_),
    .ZN(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3782_ (.I(_1565_),
    .Z(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3783_ (.I(_1532_),
    .Z(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3784_ (.A1(_2942_),
    .A2(_2943_),
    .ZN(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3785_ (.I(_1620_),
    .Z(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3786_ (.A1(_2945_),
    .A2(_2785_),
    .ZN(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3787_ (.A1(_2860_),
    .A2(_2946_),
    .ZN(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3788_ (.I(_0773_),
    .Z(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3789_ (.I(_2787_),
    .Z(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3790_ (.I(_1598_),
    .Z(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3791_ (.A1(_2948_),
    .A2(_2949_),
    .B1(_2950_),
    .B2(_1367_),
    .ZN(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3792_ (.A1(_2947_),
    .A2(_2951_),
    .Z(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3793_ (.A1(_2944_),
    .A2(_2952_),
    .ZN(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3794_ (.A1(_2941_),
    .A2(_2953_),
    .Z(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3795_ (.A1(_2929_),
    .A2(_2936_),
    .A3(_2954_),
    .ZN(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3796_ (.A1(_2888_),
    .A2(_2896_),
    .ZN(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3797_ (.A1(_2886_),
    .A2(_2897_),
    .B(_2956_),
    .ZN(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3798_ (.A1(_2825_),
    .A2(_2826_),
    .B1(_2891_),
    .B2(_2895_),
    .ZN(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3799_ (.A1(_2525_),
    .A2(_1191_),
    .ZN(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3800_ (.A1(_1224_),
    .A2(_2704_),
    .ZN(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3801_ (.I(_1158_),
    .Z(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3802_ (.A1(_2893_),
    .A2(_2961_),
    .ZN(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3803_ (.A1(_2959_),
    .A2(_2960_),
    .A3(_2962_),
    .ZN(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3804_ (.A1(_2958_),
    .A2(_2963_),
    .ZN(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3805_ (.A1(_2876_),
    .A2(_2890_),
    .Z(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3806_ (.A1(_2829_),
    .A2(_2959_),
    .B1(_2965_),
    .B2(_2889_),
    .ZN(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3807_ (.I(_2190_),
    .Z(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3808_ (.A1(_2879_),
    .A2(_2967_),
    .B1(_2430_),
    .B2(_2812_),
    .ZN(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3809_ (.I(\B[1][6] ),
    .Z(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3810_ (.A1(_2969_),
    .A2(_2813_),
    .A3(_2267_),
    .A4(_2660_),
    .Z(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3811_ (.A1(_2968_),
    .A2(_2970_),
    .ZN(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3812_ (.A1(_2966_),
    .A2(_2971_),
    .ZN(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3813_ (.A1(_2883_),
    .A2(_2972_),
    .Z(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3814_ (.A1(_2964_),
    .A2(_2973_),
    .Z(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3815_ (.A1(_2957_),
    .A2(_2974_),
    .ZN(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3816_ (.A1(_2955_),
    .A2(_2975_),
    .Z(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3817_ (.A1(_2927_),
    .A2(_2976_),
    .Z(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3818_ (.A1(_2925_),
    .A2(_2977_),
    .ZN(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3819_ (.A1(_2914_),
    .A2(_2978_),
    .Z(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3820_ (.A1(_2912_),
    .A2(_2979_),
    .Z(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3821_ (.A1(_2903_),
    .A2(_2906_),
    .B(_2980_),
    .ZN(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3822_ (.A1(_2786_),
    .A2(_0982_),
    .ZN(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3823_ (.I(_1015_),
    .Z(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3824_ (.I(\A[3][2] ),
    .Z(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3825_ (.I(_2984_),
    .Z(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3826_ (.A1(_2983_),
    .A2(_2985_),
    .ZN(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3827_ (.A1(_1796_),
    .A2(_0927_),
    .ZN(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3828_ (.I(_2786_),
    .Z(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3829_ (.I(_1015_),
    .Z(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3830_ (.A1(_2985_),
    .A2(_2988_),
    .B1(_2922_),
    .B2(_2989_),
    .ZN(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3831_ (.A1(_2982_),
    .A2(_2986_),
    .B1(_2987_),
    .B2(_2990_),
    .ZN(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3832_ (.A1(_1466_),
    .A2(_2982_),
    .A3(_0938_),
    .ZN(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3833_ (.A1(_2991_),
    .A2(_2992_),
    .ZN(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3834_ (.I(\A[3][0] ),
    .Z(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3835_ (.I(_2950_),
    .Z(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3836_ (.A1(_2994_),
    .A2(_2995_),
    .ZN(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3837_ (.A1(_0784_),
    .A2(_2996_),
    .ZN(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3838_ (.I(_2994_),
    .Z(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3839_ (.A1(_2948_),
    .A2(_2998_),
    .B1(_1807_),
    .B2(_2995_),
    .ZN(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3840_ (.A1(_2997_),
    .A2(_2999_),
    .ZN(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3841_ (.A1(_2991_),
    .A2(_2992_),
    .Z(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3842_ (.A1(_3000_),
    .A2(_3001_),
    .ZN(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3843_ (.A1(_2993_),
    .A2(_3002_),
    .ZN(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3844_ (.I(_2949_),
    .Z(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3845_ (.I(_3004_),
    .Z(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3846_ (.I(_1389_),
    .Z(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3847_ (.I(_3006_),
    .Z(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3848_ (.I(_1246_),
    .Z(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3849_ (.A1(_3008_),
    .A2(_2961_),
    .ZN(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3850_ (.A1(_1202_),
    .A2(_3009_),
    .ZN(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3851_ (.I(_3010_),
    .Z(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3852_ (.A1(_3005_),
    .A2(_3007_),
    .A3(_3011_),
    .ZN(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3853_ (.A1(_0806_),
    .A2(_1114_),
    .Z(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3854_ (.A1(_3012_),
    .A2(_3013_),
    .ZN(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3855_ (.I(_3007_),
    .Z(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3856_ (.A1(_3005_),
    .A2(_3015_),
    .A3(_3011_),
    .A4(_3013_),
    .Z(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3857_ (.A1(_3003_),
    .A2(_3014_),
    .B(_3016_),
    .ZN(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3858_ (.A1(_0762_),
    .A2(_0784_),
    .ZN(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3859_ (.A1(_0729_),
    .A2(_0795_),
    .ZN(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3860_ (.A1(_3018_),
    .A2(_3019_),
    .ZN(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3861_ (.A1(_3017_),
    .A2(_3020_),
    .Z(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3862_ (.A1(_3017_),
    .A2(_3020_),
    .ZN(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3863_ (.A1(_3021_),
    .A2(_3022_),
    .ZN(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3864_ (.I(_2998_),
    .Z(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3865_ (.I(_3024_),
    .Z(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3866_ (.A1(_2921_),
    .A2(_3025_),
    .ZN(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3867_ (.A1(_3023_),
    .A2(_3026_),
    .B(_3021_),
    .ZN(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3868_ (.A1(_1872_),
    .A2(_2774_),
    .ZN(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3869_ (.A1(_3003_),
    .A2(_3014_),
    .Z(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3870_ (.A1(_3004_),
    .A2(_3006_),
    .ZN(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3871_ (.A1(_3011_),
    .A2(_3030_),
    .Z(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3872_ (.I(_2961_),
    .Z(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3873_ (.I(_2299_),
    .Z(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3874_ (.I(_3033_),
    .Z(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3875_ (.I(_1323_),
    .Z(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3876_ (.A1(_2932_),
    .A2(_3032_),
    .B1(_3034_),
    .B2(_3035_),
    .ZN(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3877_ (.I(_2398_),
    .Z(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3878_ (.A1(_3037_),
    .A2(_2806_),
    .ZN(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3879_ (.I(_2113_),
    .Z(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3880_ (.I(_2810_),
    .Z(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3881_ (.A1(_3039_),
    .A2(_3040_),
    .ZN(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3882_ (.A1(_2931_),
    .A2(_2894_),
    .ZN(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3883_ (.I(_2070_),
    .Z(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3884_ (.I(_2201_),
    .Z(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3885_ (.I(_2113_),
    .Z(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3886_ (.A1(_3043_),
    .A2(_3040_),
    .B1(_3044_),
    .B2(_3045_),
    .ZN(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3887_ (.A1(_3038_),
    .A2(_3041_),
    .B1(_3042_),
    .B2(_3046_),
    .ZN(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3888_ (.A1(_2441_),
    .A2(_3038_),
    .A3(_2059_),
    .ZN(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3889_ (.A1(_3047_),
    .A2(_3048_),
    .ZN(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3890_ (.A1(_3047_),
    .A2(_3048_),
    .ZN(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3891_ (.A1(_3011_),
    .A2(_3036_),
    .A3(_3049_),
    .B(_3050_),
    .ZN(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3892_ (.A1(_1916_),
    .A2(_2234_),
    .Z(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3893_ (.A1(_3051_),
    .A2(_3052_),
    .ZN(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3894_ (.A1(_3051_),
    .A2(_3052_),
    .ZN(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3895_ (.A1(_3031_),
    .A2(_3053_),
    .B(_3054_),
    .ZN(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3896_ (.A1(_1905_),
    .A2(_2576_),
    .Z(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3897_ (.A1(_3055_),
    .A2(_3056_),
    .Z(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3898_ (.A1(_3055_),
    .A2(_3056_),
    .Z(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3899_ (.A1(_3029_),
    .A2(_3057_),
    .B(_3058_),
    .ZN(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3900_ (.A1(_2596_),
    .A2(_2773_),
    .ZN(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3901_ (.A1(_1862_),
    .A2(_3060_),
    .ZN(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3902_ (.A1(_3023_),
    .A2(_3026_),
    .ZN(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3903_ (.A1(_1862_),
    .A2(_3060_),
    .A3(_3059_),
    .Z(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3904_ (.A1(_3028_),
    .A2(_3059_),
    .A3(_3061_),
    .B1(_3062_),
    .B2(_3063_),
    .ZN(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3905_ (.A1(_1851_),
    .A2(_2837_),
    .Z(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3906_ (.A1(_3064_),
    .A2(_3065_),
    .Z(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3907_ (.A1(_3064_),
    .A2(_3065_),
    .Z(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3908_ (.A1(_3027_),
    .A2(_3066_),
    .B(_3067_),
    .ZN(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3909_ (.A1(_2839_),
    .A2(_2902_),
    .A3(_2904_),
    .Z(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3910_ (.A1(_3068_),
    .A2(_3069_),
    .Z(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3911_ (.A1(_0718_),
    .A2(_2939_),
    .ZN(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3912_ (.I(_2988_),
    .Z(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3913_ (.A1(_1807_),
    .A2(_3072_),
    .ZN(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3914_ (.A1(_2986_),
    .A2(_3071_),
    .A3(_3073_),
    .Z(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3915_ (.I(_2989_),
    .Z(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3916_ (.A1(_2994_),
    .A2(_3075_),
    .ZN(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3917_ (.A1(_3073_),
    .A2(_3076_),
    .Z(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3918_ (.A1(_3074_),
    .A2(_3077_),
    .ZN(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3919_ (.I(_2996_),
    .Z(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3920_ (.A1(_2984_),
    .A2(_0960_),
    .ZN(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3921_ (.I(_1576_),
    .Z(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3922_ (.A1(_3081_),
    .A2(_2989_),
    .ZN(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3923_ (.A1(_2989_),
    .A2(_2985_),
    .B1(_2988_),
    .B2(_3081_),
    .ZN(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3924_ (.A1(_3080_),
    .A2(_3082_),
    .B1(_3083_),
    .B2(_3071_),
    .ZN(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3925_ (.A1(_0894_),
    .A2(_3080_),
    .A3(_2987_),
    .ZN(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3926_ (.A1(_3084_),
    .A2(_3085_),
    .ZN(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3927_ (.A1(_3079_),
    .A2(_3086_),
    .Z(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3928_ (.A1(_3079_),
    .A2(_3086_),
    .ZN(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3929_ (.A1(_3078_),
    .A2(_3087_),
    .A3(_3088_),
    .Z(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3930_ (.I(_3089_),
    .ZN(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3931_ (.A1(_3079_),
    .A2(_3078_),
    .A3(_3086_),
    .Z(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3932_ (.I(_3091_),
    .ZN(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3933_ (.I(_3006_),
    .Z(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3934_ (.A1(_3093_),
    .A2(_2923_),
    .ZN(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3935_ (.I(_3037_),
    .Z(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3936_ (.I(_3095_),
    .Z(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3937_ (.A1(_2932_),
    .A2(_3096_),
    .ZN(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3938_ (.I(_2048_),
    .Z(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3939_ (.A1(_3008_),
    .A2(_3098_),
    .ZN(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3940_ (.A1(_3041_),
    .A2(_3099_),
    .A3(_3097_),
    .Z(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3941_ (.I(_3045_),
    .Z(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3942_ (.I(_3035_),
    .Z(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3943_ (.A1(_3101_),
    .A2(_3102_),
    .ZN(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3944_ (.A1(_3097_),
    .A2(_3100_),
    .A3(_3103_),
    .ZN(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3945_ (.A1(_2070_),
    .A2(_2026_),
    .ZN(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3946_ (.I(_2354_),
    .Z(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3947_ (.A1(_3039_),
    .A2(_3106_),
    .ZN(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3948_ (.I(_2882_),
    .Z(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3949_ (.A1(_2931_),
    .A2(_3043_),
    .B1(_3108_),
    .B2(_3045_),
    .ZN(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3950_ (.A1(_3105_),
    .A2(_3107_),
    .B1(_3109_),
    .B2(_3099_),
    .ZN(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3951_ (.A1(_2015_),
    .A2(_3105_),
    .A3(_3042_),
    .ZN(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3952_ (.A1(_3009_),
    .A2(_3110_),
    .A3(_3111_),
    .ZN(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3953_ (.A1(_3104_),
    .A2(_3112_),
    .ZN(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3954_ (.A1(_3104_),
    .A2(_3112_),
    .ZN(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3955_ (.A1(_3094_),
    .A2(_3113_),
    .B(_3114_),
    .ZN(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3956_ (.I(_2943_),
    .Z(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3957_ (.A1(_3006_),
    .A2(_3116_),
    .ZN(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3958_ (.A1(_3110_),
    .A2(_3111_),
    .ZN(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3959_ (.A1(_3110_),
    .A2(_3111_),
    .ZN(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3960_ (.A1(_3009_),
    .A2(_3118_),
    .B(_3119_),
    .ZN(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3961_ (.A1(_3010_),
    .A2(_3036_),
    .ZN(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3962_ (.A1(_3047_),
    .A2(_3048_),
    .Z(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3963_ (.A1(_3121_),
    .A2(_3122_),
    .Z(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3964_ (.A1(_3117_),
    .A2(_3120_),
    .A3(_3123_),
    .ZN(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3965_ (.A1(_3115_),
    .A2(_3124_),
    .ZN(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3966_ (.A1(_3115_),
    .A2(_3124_),
    .ZN(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3967_ (.A1(_3092_),
    .A2(_3125_),
    .B(_3126_),
    .ZN(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3968_ (.A1(_3084_),
    .A2(_3085_),
    .ZN(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3969_ (.A1(_3128_),
    .A2(_3087_),
    .ZN(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3970_ (.A1(_3000_),
    .A2(_3001_),
    .Z(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3971_ (.A1(_3129_),
    .A2(_3130_),
    .Z(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3972_ (.A1(_3120_),
    .A2(_3123_),
    .ZN(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3973_ (.A1(_3120_),
    .A2(_3123_),
    .ZN(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3974_ (.A1(_3117_),
    .A2(_3132_),
    .B(_3133_),
    .ZN(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3975_ (.A1(_3031_),
    .A2(_3053_),
    .Z(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3976_ (.A1(_3131_),
    .A2(_3134_),
    .A3(_3135_),
    .Z(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3977_ (.A1(_3127_),
    .A2(_3136_),
    .ZN(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3978_ (.A1(_3127_),
    .A2(_3136_),
    .ZN(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3979_ (.A1(_3090_),
    .A2(_3137_),
    .B(_3138_),
    .ZN(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3980_ (.A1(_3129_),
    .A2(_3130_),
    .ZN(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3981_ (.A1(_2997_),
    .A2(_3140_),
    .Z(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3982_ (.A1(_3134_),
    .A2(_3135_),
    .Z(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3983_ (.A1(_3134_),
    .A2(_3135_),
    .Z(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3984_ (.A1(_3131_),
    .A2(_3142_),
    .B(_3143_),
    .ZN(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3985_ (.A1(_3029_),
    .A2(_3057_),
    .ZN(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3986_ (.A1(_3141_),
    .A2(_3144_),
    .A3(_3145_),
    .ZN(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3987_ (.A1(_3139_),
    .A2(_3146_),
    .ZN(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3988_ (.A1(_0784_),
    .A2(_3079_),
    .A3(_3140_),
    .ZN(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3989_ (.A1(_3144_),
    .A2(_3145_),
    .Z(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3990_ (.A1(_3144_),
    .A2(_3145_),
    .Z(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3991_ (.A1(_3141_),
    .A2(_3149_),
    .B(_3150_),
    .ZN(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3992_ (.A1(_3062_),
    .A2(_3063_),
    .Z(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3993_ (.A1(_3148_),
    .A2(_3151_),
    .A3(_3152_),
    .ZN(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3994_ (.A1(_3147_),
    .A2(_3153_),
    .ZN(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3995_ (.A1(_3115_),
    .A2(_3124_),
    .A3(_3091_),
    .Z(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3996_ (.I(_3077_),
    .ZN(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3997_ (.A1(_3074_),
    .A2(_3156_),
    .Z(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3998_ (.A1(_3097_),
    .A2(_3103_),
    .ZN(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3999_ (.A1(_3100_),
    .A2(_3158_),
    .Z(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4000_ (.A1(_3093_),
    .A2(_2849_),
    .ZN(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4001_ (.A1(_3159_),
    .A2(_3160_),
    .ZN(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4002_ (.A1(_3104_),
    .A2(_3112_),
    .A3(_3094_),
    .ZN(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4003_ (.A1(_3161_),
    .A2(_3162_),
    .ZN(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4004_ (.A1(_3161_),
    .A2(_3162_),
    .ZN(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4005_ (.A1(_3157_),
    .A2(_3163_),
    .B(_3164_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4006_ (.A1(_3155_),
    .A2(_3165_),
    .ZN(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4007_ (.A1(_3161_),
    .A2(_3162_),
    .A3(_3157_),
    .ZN(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4008_ (.A1(_3100_),
    .A2(_3158_),
    .A3(_3160_),
    .Z(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4009_ (.I(_3096_),
    .Z(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4010_ (.A1(_3102_),
    .A2(_3169_),
    .ZN(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4011_ (.A1(_3015_),
    .A2(_1818_),
    .ZN(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4012_ (.A1(_3107_),
    .A2(_3170_),
    .B(_3171_),
    .C(_3158_),
    .ZN(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4013_ (.A1(_3168_),
    .A2(_3172_),
    .ZN(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4014_ (.I(_3072_),
    .Z(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4015_ (.A1(_3025_),
    .A2(_3174_),
    .ZN(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4016_ (.A1(_3082_),
    .A2(_3175_),
    .B(_3156_),
    .ZN(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4017_ (.A1(_3168_),
    .A2(_3172_),
    .Z(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4018_ (.A1(_3176_),
    .A2(_3177_),
    .ZN(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4019_ (.A1(_3173_),
    .A2(_3178_),
    .ZN(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4020_ (.A1(_3167_),
    .A2(_3179_),
    .Z(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4021_ (.I(_3093_),
    .Z(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4022_ (.I(_3181_),
    .Z(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4023_ (.A1(_3107_),
    .A2(_3170_),
    .B(_3158_),
    .ZN(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4024_ (.A1(_3182_),
    .A2(_1829_),
    .B(_3183_),
    .ZN(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4025_ (.A1(_3024_),
    .A2(_3181_),
    .ZN(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4026_ (.A1(_3103_),
    .A2(_3185_),
    .Z(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4027_ (.A1(_3183_),
    .A2(_3171_),
    .A3(_3186_),
    .ZN(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4028_ (.A1(_3076_),
    .A2(_3187_),
    .Z(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4029_ (.A1(_3172_),
    .A2(_3184_),
    .A3(_3186_),
    .B(_3188_),
    .ZN(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4030_ (.A1(_3176_),
    .A2(_3177_),
    .Z(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4031_ (.A1(_3189_),
    .A2(_3190_),
    .Z(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4032_ (.A1(_3180_),
    .A2(_3191_),
    .ZN(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4033_ (.A1(_3166_),
    .A2(_3192_),
    .Z(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4034_ (.A1(_3090_),
    .A2(_3127_),
    .A3(_3136_),
    .Z(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4035_ (.A1(_3167_),
    .A2(_3179_),
    .ZN(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4036_ (.A1(_3155_),
    .A2(_3165_),
    .ZN(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4037_ (.A1(_3166_),
    .A2(_3195_),
    .B(_3196_),
    .ZN(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4038_ (.A1(_3194_),
    .A2(_3197_),
    .Z(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4039_ (.A1(_3193_),
    .A2(_3198_),
    .Z(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4040_ (.A1(_3166_),
    .A2(_3195_),
    .A3(_3194_),
    .Z(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4041_ (.A1(_3199_),
    .A2(_3200_),
    .Z(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4042_ (.A1(_3139_),
    .A2(_3146_),
    .Z(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4043_ (.A1(_3196_),
    .A2(_3194_),
    .ZN(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4044_ (.A1(_3202_),
    .A2(_3203_),
    .ZN(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4045_ (.A1(_3201_),
    .A2(_3204_),
    .ZN(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4046_ (.A1(_3202_),
    .A2(_3203_),
    .ZN(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4047_ (.A1(_3147_),
    .A2(_3206_),
    .ZN(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4048_ (.A1(_3151_),
    .A2(_3152_),
    .Z(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4049_ (.A1(_3148_),
    .A2(_3208_),
    .Z(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4050_ (.A1(_3154_),
    .A2(_3205_),
    .B1(_3207_),
    .B2(_3209_),
    .ZN(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4051_ (.A1(_3027_),
    .A2(_3066_),
    .ZN(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4052_ (.A1(_3151_),
    .A2(_3152_),
    .Z(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4053_ (.A1(_3148_),
    .A2(_3208_),
    .B(_3212_),
    .ZN(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4054_ (.A1(_3211_),
    .A2(_3213_),
    .ZN(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4055_ (.A1(_3070_),
    .A2(_3210_),
    .A3(_3214_),
    .ZN(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4056_ (.A1(_2904_),
    .A2(_2905_),
    .ZN(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4057_ (.A1(_3027_),
    .A2(_3066_),
    .B(_3069_),
    .C(_3067_),
    .ZN(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _4058_ (.A1(_2906_),
    .A2(_3068_),
    .A3(_3216_),
    .B1(_3217_),
    .B2(_3211_),
    .B3(_3213_),
    .ZN(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4059_ (.A1(_2904_),
    .A2(_2905_),
    .B(_2903_),
    .ZN(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4060_ (.A1(_2980_),
    .A2(_3219_),
    .ZN(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4061_ (.A1(_3215_),
    .A2(_3218_),
    .B(_3220_),
    .ZN(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4062_ (.A1(_2981_),
    .A2(_3221_),
    .ZN(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4063_ (.A1(_2914_),
    .A2(_2978_),
    .ZN(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4064_ (.A1(_2912_),
    .A2(_2979_),
    .B(_3223_),
    .ZN(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4065_ (.I(_2923_),
    .Z(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4066_ (.A1(_2908_),
    .A2(_3225_),
    .A3(_2920_),
    .ZN(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4067_ (.A1(_2916_),
    .A2(_2919_),
    .B(_3226_),
    .ZN(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4068_ (.I(_3227_),
    .ZN(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4069_ (.A1(_2927_),
    .A2(_2976_),
    .ZN(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4070_ (.A1(_2925_),
    .A2(_2977_),
    .ZN(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4071_ (.A1(_3229_),
    .A2(_3230_),
    .ZN(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4072_ (.A1(_2907_),
    .A2(_3116_),
    .ZN(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4073_ (.A1(_2944_),
    .A2(_2952_),
    .ZN(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4074_ (.A1(_2947_),
    .A2(_3233_),
    .ZN(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4075_ (.A1(_2936_),
    .A2(_2954_),
    .Z(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4076_ (.A1(_2936_),
    .A2(_2954_),
    .Z(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4077_ (.A1(_2929_),
    .A2(_3235_),
    .B(_3236_),
    .ZN(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4078_ (.A1(_3234_),
    .A2(_3237_),
    .Z(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4079_ (.A1(_3232_),
    .A2(_3238_),
    .Z(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4080_ (.A1(_2957_),
    .A2(_2974_),
    .ZN(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4081_ (.A1(_2955_),
    .A2(_2975_),
    .B(_3240_),
    .ZN(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4082_ (.A1(_2867_),
    .A2(_2868_),
    .B1(_2941_),
    .B2(_2953_),
    .ZN(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4083_ (.I(_2930_),
    .Z(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4084_ (.I(_2879_),
    .Z(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4085_ (.I(_3244_),
    .Z(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4086_ (.I(_3108_),
    .Z(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4087_ (.I(_3044_),
    .Z(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4088_ (.A1(_3243_),
    .A2(_3245_),
    .A3(_3246_),
    .A4(_3247_),
    .ZN(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4089_ (.A1(_2966_),
    .A2(_2971_),
    .ZN(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4090_ (.A1(_3248_),
    .A2(_2972_),
    .B(_3249_),
    .ZN(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4091_ (.I(_0707_),
    .Z(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4092_ (.A1(_3251_),
    .A2(_2949_),
    .ZN(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4093_ (.A1(_2937_),
    .A2(_2950_),
    .ZN(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4094_ (.A1(_2946_),
    .A2(_3253_),
    .ZN(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4095_ (.A1(_3252_),
    .A2(_3254_),
    .Z(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4096_ (.A1(_3250_),
    .A2(_3255_),
    .Z(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4097_ (.A1(_3242_),
    .A2(_3256_),
    .ZN(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4098_ (.A1(_2958_),
    .A2(_2963_),
    .ZN(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4099_ (.A1(_2964_),
    .A2(_2973_),
    .B(_3258_),
    .ZN(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4100_ (.I(_2892_),
    .Z(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4101_ (.A1(_3260_),
    .A2(_3034_),
    .ZN(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4102_ (.I(_2343_),
    .Z(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4103_ (.I(_2821_),
    .Z(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4104_ (.I(_3263_),
    .Z(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4105_ (.A1(_3262_),
    .A2(_3264_),
    .ZN(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4106_ (.A1(_3260_),
    .A2(_1235_),
    .ZN(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4107_ (.A1(_2959_),
    .A2(_3266_),
    .ZN(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4108_ (.A1(_3261_),
    .A2(_3265_),
    .B(_3267_),
    .ZN(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4109_ (.I(_2704_),
    .Z(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4110_ (.I(_3269_),
    .Z(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4111_ (.I(_2081_),
    .Z(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4112_ (.I(_3271_),
    .Z(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4113_ (.A1(_1312_),
    .A2(_3270_),
    .B1(_3244_),
    .B2(_3272_),
    .ZN(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4114_ (.I(_2969_),
    .Z(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4115_ (.A1(_3274_),
    .A2(_3269_),
    .A3(_3244_),
    .A4(_3271_),
    .Z(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4116_ (.A1(_3273_),
    .A2(_3275_),
    .ZN(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4117_ (.A1(_2959_),
    .A2(_2962_),
    .Z(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4118_ (.A1(_2890_),
    .A2(_3261_),
    .B1(_3277_),
    .B2(_2960_),
    .ZN(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4119_ (.A1(_3276_),
    .A2(_3278_),
    .Z(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4120_ (.A1(_2970_),
    .A2(_3279_),
    .Z(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4121_ (.A1(_3268_),
    .A2(_3280_),
    .Z(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4122_ (.A1(_3259_),
    .A2(_3281_),
    .ZN(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4123_ (.A1(_3257_),
    .A2(_3282_),
    .Z(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4124_ (.A1(_3241_),
    .A2(_3283_),
    .ZN(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4125_ (.A1(_3239_),
    .A2(_3284_),
    .Z(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4126_ (.A1(_3228_),
    .A2(_3231_),
    .A3(_3285_),
    .Z(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4127_ (.A1(_3224_),
    .A2(_3286_),
    .Z(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4128_ (.I(net16),
    .ZN(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4129_ (.I(net15),
    .ZN(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4130_ (.A1(_3288_),
    .A2(_3289_),
    .ZN(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4131_ (.I(_3290_),
    .Z(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4132_ (.A1(_3222_),
    .A2(_3287_),
    .B(_3291_),
    .ZN(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4133_ (.A1(_3222_),
    .A2(_3287_),
    .B(_3292_),
    .ZN(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4134_ (.A1(_0696_),
    .A2(_3293_),
    .ZN(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4135_ (.I(_3288_),
    .Z(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4136_ (.I(_3295_),
    .Z(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4137_ (.I(\A[1][0] ),
    .Z(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4138_ (.A1(_2942_),
    .A2(_3297_),
    .ZN(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4139_ (.I(\A[1][2] ),
    .Z(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4140_ (.A1(_3299_),
    .A2(_0751_),
    .ZN(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4141_ (.I(\A[1][1] ),
    .Z(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4142_ (.A1(_2945_),
    .A2(_3301_),
    .ZN(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4143_ (.A1(_3300_),
    .A2(_3302_),
    .ZN(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4144_ (.A1(_3298_),
    .A2(_3303_),
    .ZN(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4145_ (.I(\A[1][4] ),
    .Z(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4146_ (.A1(_2863_),
    .A2(_3305_),
    .ZN(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4147_ (.I(_0861_),
    .Z(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4148_ (.I(\A[1][3] ),
    .Z(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4149_ (.I(_3308_),
    .Z(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4150_ (.A1(_3307_),
    .A2(_3309_),
    .ZN(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4151_ (.I(_3299_),
    .Z(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4152_ (.A1(_3311_),
    .A2(_0927_),
    .ZN(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4153_ (.I(_3305_),
    .Z(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4154_ (.A1(_0971_),
    .A2(_3309_),
    .B1(_3313_),
    .B2(_3307_),
    .ZN(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4155_ (.A1(_3306_),
    .A2(_3310_),
    .B1(_3312_),
    .B2(_3314_),
    .ZN(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4156_ (.A1(\A[1][5] ),
    .A2(_1510_),
    .ZN(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4157_ (.I(\A[1][3] ),
    .Z(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4158_ (.A1(_3317_),
    .A2(_0927_),
    .ZN(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4159_ (.A1(_3306_),
    .A2(_3316_),
    .A3(_3318_),
    .ZN(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4160_ (.A1(_3315_),
    .A2(_3319_),
    .ZN(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4161_ (.A1(_3315_),
    .A2(_3319_),
    .ZN(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4162_ (.A1(_3304_),
    .A2(_3320_),
    .B(_3321_),
    .ZN(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4163_ (.I(\A[0][2] ),
    .Z(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4164_ (.A1(_3323_),
    .A2(_2651_),
    .ZN(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4165_ (.I(\A[0][1] ),
    .Z(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4166_ (.A1(_3325_),
    .A2(_2310_),
    .ZN(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4167_ (.A1(_3324_),
    .A2(_3326_),
    .ZN(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4168_ (.I(\A[0][0] ),
    .Z(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4169_ (.A1(_3262_),
    .A2(_3328_),
    .ZN(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4170_ (.A1(_3324_),
    .A2(_3326_),
    .ZN(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4171_ (.A1(_3329_),
    .A2(_3330_),
    .ZN(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4172_ (.A1(_1312_),
    .A2(_3328_),
    .ZN(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4173_ (.I(\A[1][6] ),
    .Z(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4174_ (.I(_3333_),
    .Z(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4175_ (.A1(_3334_),
    .A2(_1389_),
    .ZN(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4176_ (.A1(_3332_),
    .A2(_3335_),
    .Z(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4177_ (.A1(_3332_),
    .A2(_3335_),
    .ZN(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4178_ (.A1(_3327_),
    .A2(_3331_),
    .B(_3336_),
    .C(_3337_),
    .ZN(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4179_ (.A1(_0707_),
    .A2(_3301_),
    .ZN(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4180_ (.A1(_0773_),
    .A2(\A[1][2] ),
    .ZN(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4181_ (.A1(\A[1][3] ),
    .A2(_1598_),
    .ZN(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4182_ (.A1(_3340_),
    .A2(_3341_),
    .ZN(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4183_ (.A1(_3339_),
    .A2(_3342_),
    .ZN(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4184_ (.A1(_3307_),
    .A2(_3313_),
    .ZN(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4185_ (.I(\A[1][5] ),
    .Z(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4186_ (.I(_3345_),
    .Z(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4187_ (.A1(_3346_),
    .A2(_2786_),
    .ZN(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4188_ (.A1(_3306_),
    .A2(_3316_),
    .Z(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4189_ (.A1(_3344_),
    .A2(_3347_),
    .B1(_3348_),
    .B2(_3318_),
    .ZN(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4190_ (.I(\A[1][6] ),
    .Z(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4191_ (.I(_3350_),
    .Z(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4192_ (.A1(_3351_),
    .A2(_1015_),
    .ZN(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4193_ (.I(_3305_),
    .Z(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4194_ (.A1(_2939_),
    .A2(_3353_),
    .ZN(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4195_ (.A1(_3347_),
    .A2(_3352_),
    .A3(_3354_),
    .ZN(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4196_ (.A1(_3343_),
    .A2(_3349_),
    .A3(_3355_),
    .Z(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4197_ (.A1(_3338_),
    .A2(_3356_),
    .Z(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4198_ (.A1(_3338_),
    .A2(_3356_),
    .ZN(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4199_ (.A1(_3322_),
    .A2(_3357_),
    .B(_3358_),
    .ZN(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4200_ (.A1(_2945_),
    .A2(_3317_),
    .ZN(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4201_ (.A1(_3300_),
    .A2(_3360_),
    .ZN(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4202_ (.A1(_3339_),
    .A2(_3342_),
    .ZN(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4203_ (.A1(_3361_),
    .A2(_3362_),
    .ZN(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4204_ (.A1(_3359_),
    .A2(_3363_),
    .Z(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4205_ (.A1(_3359_),
    .A2(_3363_),
    .ZN(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4206_ (.A1(_3364_),
    .A2(_3365_),
    .ZN(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4207_ (.I(_3301_),
    .Z(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4208_ (.I(_3367_),
    .Z(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4209_ (.I(_3368_),
    .Z(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4210_ (.A1(_2921_),
    .A2(_3369_),
    .ZN(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4211_ (.A1(_3366_),
    .A2(_3370_),
    .B(_3364_),
    .ZN(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4212_ (.A1(_3366_),
    .A2(_3370_),
    .Z(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4213_ (.A1(_3322_),
    .A2(_3357_),
    .Z(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4214_ (.I(_3373_),
    .ZN(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4215_ (.A1(_3327_),
    .A2(_3331_),
    .ZN(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4216_ (.A1(_3336_),
    .A2(_3337_),
    .ZN(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4217_ (.A1(_3375_),
    .A2(_3376_),
    .ZN(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4218_ (.A1(_3329_),
    .A2(_3330_),
    .ZN(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4219_ (.I(\A[0][4] ),
    .Z(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4220_ (.I(_3379_),
    .Z(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4221_ (.A1(_3037_),
    .A2(_3380_),
    .ZN(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4222_ (.I(\A[0][3] ),
    .Z(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4223_ (.I(_3382_),
    .Z(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4224_ (.A1(_3045_),
    .A2(_3383_),
    .ZN(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4225_ (.I(_3323_),
    .Z(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4226_ (.A1(_3385_),
    .A2(_2894_),
    .ZN(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4227_ (.I(_3380_),
    .Z(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4228_ (.A1(_3095_),
    .A2(_3383_),
    .B1(_3387_),
    .B2(_1982_),
    .ZN(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4229_ (.A1(_3381_),
    .A2(_3384_),
    .B1(_3386_),
    .B2(_3388_),
    .ZN(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4230_ (.I(\A[0][3] ),
    .Z(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4231_ (.A1(_2048_),
    .A2(_3390_),
    .ZN(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4232_ (.I(\A[0][5] ),
    .Z(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4233_ (.I(_3392_),
    .Z(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4234_ (.A1(_3393_),
    .A2(_2419_),
    .ZN(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4235_ (.A1(_3381_),
    .A2(_3391_),
    .A3(_3394_),
    .ZN(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4236_ (.A1(_3389_),
    .A2(_3395_),
    .ZN(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4237_ (.A1(_3389_),
    .A2(_3395_),
    .ZN(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4238_ (.A1(_3378_),
    .A2(_3396_),
    .B(_3397_),
    .ZN(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4239_ (.I(\A[0][2] ),
    .Z(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4240_ (.A1(_3399_),
    .A2(_2310_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4241_ (.I(_3325_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4242_ (.A1(_2343_),
    .A2(_0065_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4243_ (.A1(_3382_),
    .A2(_1158_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4244_ (.A1(_0064_),
    .A2(_0066_),
    .A3(_0067_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4245_ (.I(_3379_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4246_ (.I(_0069_),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4247_ (.A1(_1982_),
    .A2(_0070_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4248_ (.I(\A[0][5] ),
    .Z(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4249_ (.I(_0072_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4250_ (.A1(_0073_),
    .A2(_2697_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4251_ (.I(_3393_),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4252_ (.A1(_0075_),
    .A2(_1982_),
    .B1(_3095_),
    .B2(_3387_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4253_ (.A1(_0071_),
    .A2(_0074_),
    .B1(_0076_),
    .B2(_3391_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4254_ (.A1(_2037_),
    .A2(_0069_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4255_ (.I(\A[0][6] ),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4256_ (.I(_0079_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4257_ (.A1(_0080_),
    .A2(_2113_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4258_ (.A1(_0074_),
    .A2(_0078_),
    .A3(_0081_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4259_ (.A1(_0077_),
    .A2(_0082_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4260_ (.A1(_0068_),
    .A2(_0083_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4261_ (.A1(_3398_),
    .A2(_0084_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4262_ (.A1(_3398_),
    .A2(_0084_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4263_ (.A1(_3377_),
    .A2(_0085_),
    .B(_0086_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4264_ (.I(\A[0][3] ),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4265_ (.A1(_0088_),
    .A2(_3033_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4266_ (.A1(_0064_),
    .A2(_0067_),
    .Z(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4267_ (.A1(_3324_),
    .A2(_0089_),
    .B1(_0090_),
    .B2(_0066_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4268_ (.A1(\A[1][7] ),
    .A2(\B[3][0] ),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4269_ (.A1(\B[1][6] ),
    .A2(_2765_),
    .A3(\A[0][0] ),
    .A4(\A[0][1] ),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4270_ (.A1(_2763_),
    .A2(\A[0][0] ),
    .B1(\A[0][1] ),
    .B2(_2762_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4271_ (.A1(_0092_),
    .A2(_0093_),
    .A3(_0094_),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4272_ (.A1(_0093_),
    .A2(_0094_),
    .B(_0092_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4273_ (.A1(_0095_),
    .A2(_0096_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4274_ (.A1(_0091_),
    .A2(_0097_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4275_ (.A1(_3336_),
    .A2(_0098_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4276_ (.A1(_0077_),
    .A2(_0082_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4277_ (.A1(_0068_),
    .A2(_0083_),
    .B(_0100_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4278_ (.I(\A[0][6] ),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4279_ (.A1(_0102_),
    .A2(_2398_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4280_ (.A1(_0080_),
    .A2(_2419_),
    .B1(_3037_),
    .B2(_3393_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4281_ (.A1(_3394_),
    .A2(_0103_),
    .B1(_0104_),
    .B2(_0078_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4282_ (.A1(_0072_),
    .A2(_2484_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4283_ (.I(\A[0][7] ),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4284_ (.A1(_0107_),
    .A2(_1971_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4285_ (.A1(_0103_),
    .A2(_0106_),
    .A3(_0108_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4286_ (.A1(_0105_),
    .A2(_0109_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4287_ (.I(\A[0][4] ),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4288_ (.I(_0111_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4289_ (.A1(_2651_),
    .A2(_0112_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4290_ (.I(_3399_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4291_ (.A1(_1235_),
    .A2(_0114_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4292_ (.A1(_0089_),
    .A2(_0113_),
    .A3(_0115_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4293_ (.A1(_0110_),
    .A2(_0116_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4294_ (.A1(_0099_),
    .A2(_0101_),
    .A3(_0117_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4295_ (.A1(_0087_),
    .A2(_0118_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4296_ (.A1(_0087_),
    .A2(_0118_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4297_ (.A1(_3374_),
    .A2(_0119_),
    .B(_0120_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4298_ (.A1(_3349_),
    .A2(_3355_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4299_ (.A1(_3349_),
    .A2(_3355_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4300_ (.A1(_3343_),
    .A2(_0122_),
    .B(_0123_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4301_ (.A1(_0091_),
    .A2(_0097_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4302_ (.A1(_3336_),
    .A2(_0098_),
    .B(_0125_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4303_ (.A1(_3251_),
    .A2(_3311_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4304_ (.I(\A[1][4] ),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4305_ (.A1(_0128_),
    .A2(_0751_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4306_ (.A1(_3360_),
    .A2(_0129_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4307_ (.A1(_0127_),
    .A2(_0130_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4308_ (.A1(_3350_),
    .A2(_2863_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4309_ (.I(_3345_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4310_ (.A1(_3351_),
    .A2(_3307_),
    .B1(_2988_),
    .B2(_0133_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4311_ (.A1(_3316_),
    .A2(_0132_),
    .B1(_0134_),
    .B2(_3354_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4312_ (.I(\A[1][7] ),
    .Z(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4313_ (.A1(_0136_),
    .A2(_1004_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4314_ (.A1(_3345_),
    .A2(_1081_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4315_ (.A1(_0132_),
    .A2(_0137_),
    .A3(_0138_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4316_ (.A1(_0135_),
    .A2(_0139_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4317_ (.A1(_0131_),
    .A2(_0140_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4318_ (.A1(_0124_),
    .A2(_0126_),
    .A3(_0141_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4319_ (.A1(_0101_),
    .A2(_0117_),
    .ZN(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4320_ (.A1(_0101_),
    .A2(_0117_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4321_ (.A1(_0099_),
    .A2(_0143_),
    .B(_0144_),
    .ZN(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4322_ (.A1(_0092_),
    .A2(_0093_),
    .A3(_0094_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4323_ (.A1(_0093_),
    .A2(_0146_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4324_ (.A1(_0111_),
    .A2(_1191_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4325_ (.I(_3382_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4326_ (.A1(_2961_),
    .A2(_0070_),
    .B1(_3033_),
    .B2(_0149_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4327_ (.A1(_0067_),
    .A2(_0148_),
    .B1(_0150_),
    .B2(_0115_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4328_ (.I(_3325_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4329_ (.A1(_2809_),
    .A2(_0152_),
    .B1(_3385_),
    .B2(_3274_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4330_ (.A1(_3274_),
    .A2(_2809_),
    .A3(_0152_),
    .A4(_0114_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4331_ (.A1(_0153_),
    .A2(_0154_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4332_ (.A1(_0151_),
    .A2(_0155_),
    .Z(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4333_ (.A1(_0147_),
    .A2(_0156_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4334_ (.A1(_0105_),
    .A2(_0109_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4335_ (.A1(_0110_),
    .A2(_0116_),
    .B(_0158_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4336_ (.A1(_3392_),
    .A2(_2644_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4337_ (.I(\A[0][3] ),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4338_ (.A1(_2343_),
    .A2(_0161_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4339_ (.A1(_0148_),
    .A2(_0160_),
    .A3(_0162_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4340_ (.I(\A[0][7] ),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4341_ (.A1(_0164_),
    .A2(_1938_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4342_ (.A1(_0102_),
    .A2(_2037_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4343_ (.A1(_0165_),
    .A2(_0166_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4344_ (.I(\A[0][6] ),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4345_ (.A1(_0107_),
    .A2(_1971_),
    .B1(_2697_),
    .B2(_0168_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4346_ (.A1(_0107_),
    .A2(_0079_),
    .A3(_2102_),
    .A4(_2697_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4347_ (.A1(_0106_),
    .A2(_0169_),
    .B(_0170_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4348_ (.A1(_0167_),
    .A2(_0171_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4349_ (.A1(_0163_),
    .A2(_0172_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4350_ (.A1(_0159_),
    .A2(_0173_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4351_ (.A1(_0157_),
    .A2(_0174_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4352_ (.A1(_0145_),
    .A2(_0175_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4353_ (.A1(_0142_),
    .A2(_0176_),
    .Z(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4354_ (.A1(_0121_),
    .A2(_0177_),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4355_ (.A1(_0121_),
    .A2(_0177_),
    .Z(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4356_ (.A1(_3372_),
    .A2(_0178_),
    .B(_0179_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4357_ (.A1(_0126_),
    .A2(_0141_),
    .Z(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4358_ (.A1(_0126_),
    .A2(_0141_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4359_ (.A1(_0124_),
    .A2(_0181_),
    .B(_0182_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4360_ (.A1(_1620_),
    .A2(\A[1][4] ),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4361_ (.A1(_3341_),
    .A2(_0184_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4362_ (.A1(_0127_),
    .A2(_0130_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4363_ (.A1(_0185_),
    .A2(_0186_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4364_ (.A1(_0183_),
    .A2(_0187_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4365_ (.I(_3311_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4366_ (.I(_0189_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4367_ (.I(_0190_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4368_ (.A1(_2921_),
    .A2(_0191_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4369_ (.A1(_0188_),
    .A2(_0192_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4370_ (.A1(_0145_),
    .A2(_0175_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4371_ (.A1(_0142_),
    .A2(_0176_),
    .B(_0194_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4372_ (.A1(_0131_),
    .A2(_0140_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4373_ (.A1(_0135_),
    .A2(_0139_),
    .B(_0196_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4374_ (.A1(_0151_),
    .A2(_0155_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4375_ (.A1(_0151_),
    .A2(_0155_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4376_ (.A1(_0147_),
    .A2(_0198_),
    .B(_0199_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4377_ (.A1(_1565_),
    .A2(_3308_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4378_ (.A1(\A[1][5] ),
    .A2(\B[3][4] ),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4379_ (.A1(_0184_),
    .A2(_0202_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4380_ (.A1(_0201_),
    .A2(_0203_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4381_ (.A1(_0136_),
    .A2(_1004_),
    .B1(_0960_),
    .B2(_3350_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4382_ (.A1(_0136_),
    .A2(_3333_),
    .A3(_1004_),
    .A4(_0960_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4383_ (.A1(_0205_),
    .A2(_0138_),
    .B(_0206_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4384_ (.A1(\A[1][7] ),
    .A2(_0817_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4385_ (.A1(\A[1][6] ),
    .A2(_0916_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4386_ (.A1(_0208_),
    .A2(_0209_),
    .Z(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4387_ (.A1(_0207_),
    .A2(_0210_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4388_ (.A1(_0204_),
    .A2(_0211_),
    .Z(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4389_ (.A1(_0200_),
    .A2(_0212_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4390_ (.A1(_0197_),
    .A2(_0213_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4391_ (.A1(_0159_),
    .A2(_0173_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4392_ (.A1(_0157_),
    .A2(_0174_),
    .B(_0215_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4393_ (.A1(_0072_),
    .A2(\B[1][4] ),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4394_ (.A1(_0148_),
    .A2(_0160_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4395_ (.A1(_0113_),
    .A2(_0217_),
    .B1(_0218_),
    .B2(_0162_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4396_ (.I(_3399_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4397_ (.A1(_2879_),
    .A2(_0220_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4398_ (.A1(_1301_),
    .A2(_0088_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4399_ (.A1(_2969_),
    .A2(_2813_),
    .A3(_3323_),
    .A4(_0161_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4400_ (.A1(_0221_),
    .A2(_0222_),
    .B(_0223_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4401_ (.A1(_0219_),
    .A2(_0224_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4402_ (.A1(_0154_),
    .A2(_0225_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4403_ (.A1(_0167_),
    .A2(_0171_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4404_ (.A1(_0163_),
    .A2(_0172_),
    .B(_0227_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4405_ (.I(_0164_),
    .Z(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4406_ (.I(_0229_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4407_ (.A1(_0230_),
    .A2(_2894_),
    .A3(_0103_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4408_ (.A1(_2332_),
    .A2(_3379_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4409_ (.A1(_0102_),
    .A2(\B[1][3] ),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4410_ (.A1(_0217_),
    .A2(_0232_),
    .A3(_0233_),
    .Z(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4411_ (.A1(_0231_),
    .A2(_0234_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4412_ (.A1(_0228_),
    .A2(_0235_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4413_ (.A1(_0226_),
    .A2(_0236_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4414_ (.A1(_0216_),
    .A2(_0237_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4415_ (.A1(_0214_),
    .A2(_0238_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4416_ (.A1(_0195_),
    .A2(_0239_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4417_ (.A1(_0193_),
    .A2(_0240_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4418_ (.A1(_0180_),
    .A2(_0241_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4419_ (.A1(_0180_),
    .A2(_0241_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4420_ (.A1(_3371_),
    .A2(_0242_),
    .B(_0243_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4421_ (.A1(_0183_),
    .A2(_0187_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4422_ (.A1(_0188_),
    .A2(_0192_),
    .B(_0245_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4423_ (.A1(_0195_),
    .A2(_0239_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4424_ (.A1(_0193_),
    .A2(_0240_),
    .B(_0247_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4425_ (.A1(_0197_),
    .A2(_0213_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4426_ (.A1(_0200_),
    .A2(_0212_),
    .B(_0249_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4427_ (.A1(_0184_),
    .A2(_0202_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4428_ (.A1(_0201_),
    .A2(_0203_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4429_ (.A1(_0251_),
    .A2(_0252_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4430_ (.A1(_0250_),
    .A2(_0253_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4431_ (.I(_3308_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4432_ (.I(_0255_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4433_ (.I(_0256_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4434_ (.A1(_1785_),
    .A2(_0257_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4435_ (.A1(_0254_),
    .A2(_0258_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4436_ (.A1(_0216_),
    .A2(_0237_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4437_ (.A1(_0214_),
    .A2(_0238_),
    .B(_0260_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4438_ (.A1(_0228_),
    .A2(_0235_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4439_ (.A1(_0226_),
    .A2(_0236_),
    .B(_0262_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4440_ (.A1(_0165_),
    .A2(_0166_),
    .B1(_0231_),
    .B2(_0234_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4441_ (.A1(_0079_),
    .A2(_2299_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4442_ (.A1(_3392_),
    .A2(_2332_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4443_ (.A1(_0107_),
    .A2(_2644_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4444_ (.A1(_0265_),
    .A2(_0266_),
    .A3(_0267_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4445_ (.A1(_0264_),
    .A2(_0268_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4446_ (.A1(_0217_),
    .A2(_0233_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4447_ (.A1(_0160_),
    .A2(_0265_),
    .B1(_0270_),
    .B2(_0232_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4448_ (.A1(_2766_),
    .A2(_3382_),
    .B1(_0069_),
    .B2(_1290_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4449_ (.A1(_2762_),
    .A2(_2763_),
    .A3(_3390_),
    .A4(_0111_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4450_ (.A1(_0272_),
    .A2(_0273_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4451_ (.A1(_0271_),
    .A2(_0274_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4452_ (.A1(_0223_),
    .A2(_0275_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4453_ (.A1(_0269_),
    .A2(_0276_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4454_ (.A1(_0263_),
    .A2(_0277_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4455_ (.A1(_0207_),
    .A2(_0210_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4456_ (.A1(_0204_),
    .A2(_0211_),
    .B(_0279_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4457_ (.I(_0065_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4458_ (.I(_0281_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4459_ (.A1(_2930_),
    .A2(_0282_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4460_ (.A1(_0219_),
    .A2(_0224_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4461_ (.A1(_0283_),
    .A2(_0221_),
    .A3(_0225_),
    .B(_0284_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4462_ (.I(\A[1][7] ),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4463_ (.I(_0286_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4464_ (.A1(_0287_),
    .A2(_2940_),
    .A3(_0132_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4465_ (.A1(_2942_),
    .A2(_3353_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4466_ (.A1(_3333_),
    .A2(_0773_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4467_ (.A1(_0202_),
    .A2(_0290_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4468_ (.A1(_3346_),
    .A2(_2945_),
    .B1(_2950_),
    .B2(_3351_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4469_ (.A1(_0291_),
    .A2(_0292_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4470_ (.A1(_0289_),
    .A2(_0293_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4471_ (.A1(_0288_),
    .A2(_0294_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4472_ (.A1(_0280_),
    .A2(_0285_),
    .A3(_0295_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4473_ (.A1(_0278_),
    .A2(_0296_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4474_ (.A1(_0261_),
    .A2(_0297_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4475_ (.A1(_0259_),
    .A2(_0298_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4476_ (.A1(_0248_),
    .A2(_0299_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4477_ (.A1(_0246_),
    .A2(_0300_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4478_ (.A1(_0244_),
    .A2(_0301_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4479_ (.I(_0302_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4480_ (.I(_0303_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4481_ (.A1(_0971_),
    .A2(_3309_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4482_ (.A1(_3075_),
    .A2(_0189_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4483_ (.I(_3301_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4484_ (.A1(_0307_),
    .A2(_2939_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4485_ (.A1(_0189_),
    .A2(_3072_),
    .B1(_0256_),
    .B2(_2983_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4486_ (.A1(_0305_),
    .A2(_0306_),
    .B1(_0308_),
    .B2(_0309_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4487_ (.A1(_3344_),
    .A2(_0305_),
    .A3(_3312_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4488_ (.A1(_0310_),
    .A2(_0311_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4489_ (.I(_3297_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4490_ (.I(_0307_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4491_ (.A1(_2948_),
    .A2(_0313_),
    .A3(_0314_),
    .A4(_2995_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4492_ (.I(_0315_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4493_ (.I(_2948_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4494_ (.I(_0313_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4495_ (.I(_2995_),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4496_ (.A1(_0317_),
    .A2(_0318_),
    .B1(_3368_),
    .B2(_0319_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4497_ (.A1(_0316_),
    .A2(_0320_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4498_ (.A1(_0310_),
    .A2(_0311_),
    .Z(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4499_ (.A1(_0321_),
    .A2(_0322_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4500_ (.A1(_0312_),
    .A2(_0323_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4501_ (.I(_0133_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4502_ (.I(_0325_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4503_ (.I(\A[0][0] ),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4504_ (.I(_0327_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4505_ (.A1(_0328_),
    .A2(_3032_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4506_ (.A1(_3326_),
    .A2(_0329_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4507_ (.I(_0330_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4508_ (.A1(_0326_),
    .A2(_3093_),
    .A3(_0331_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4509_ (.A1(_3304_),
    .A2(_3320_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4510_ (.A1(_0332_),
    .A2(_0333_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4511_ (.A1(_0326_),
    .A2(_3015_),
    .A3(_0331_),
    .A4(_0333_),
    .Z(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4512_ (.A1(_0324_),
    .A2(_0334_),
    .B(_0335_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4513_ (.A1(_3300_),
    .A2(_3302_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4514_ (.A1(_3298_),
    .A2(_3303_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4515_ (.A1(_0337_),
    .A2(_0338_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4516_ (.A1(_0336_),
    .A2(_0339_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4517_ (.I(_0318_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4518_ (.I(_0341_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4519_ (.A1(_2907_),
    .A2(_0342_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4520_ (.A1(_0336_),
    .A2(_0339_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4521_ (.A1(_0340_),
    .A2(_0343_),
    .B(_0344_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4522_ (.A1(_3374_),
    .A2(_0119_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4523_ (.A1(_0324_),
    .A2(_0334_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4524_ (.A1(_0325_),
    .A2(_3007_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4525_ (.A1(_0331_),
    .A2(_0348_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4526_ (.I(_0282_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4527_ (.I(_0328_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4528_ (.A1(_0350_),
    .A2(_3032_),
    .B1(_3034_),
    .B2(_0351_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4529_ (.A1(_3095_),
    .A2(_3383_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4530_ (.I(_3385_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4531_ (.A1(_3101_),
    .A2(_0354_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4532_ (.A1(_0281_),
    .A2(_3098_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4533_ (.I(_0149_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4534_ (.A1(_3096_),
    .A2(_0354_),
    .B1(_0357_),
    .B2(_3039_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4535_ (.A1(_0353_),
    .A2(_0355_),
    .B1(_0356_),
    .B2(_0358_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4536_ (.A1(_0071_),
    .A2(_0353_),
    .A3(_3386_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4537_ (.A1(_0359_),
    .A2(_0360_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4538_ (.A1(_0359_),
    .A2(_0360_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4539_ (.A1(_0331_),
    .A2(_0352_),
    .A3(_0361_),
    .B(_0362_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4540_ (.A1(_3378_),
    .A2(_3396_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4541_ (.A1(_0363_),
    .A2(_0364_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4542_ (.A1(_0363_),
    .A2(_0364_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4543_ (.A1(_0349_),
    .A2(_0365_),
    .B(_0366_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4544_ (.A1(_3398_),
    .A2(_0084_),
    .A3(_3377_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4545_ (.A1(_0367_),
    .A2(_0368_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4546_ (.A1(_0367_),
    .A2(_0368_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4547_ (.A1(_0347_),
    .A2(_0369_),
    .B(_0370_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4548_ (.A1(_0087_),
    .A2(_0118_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4549_ (.A1(_3373_),
    .A2(_0372_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4550_ (.A1(_0340_),
    .A2(_0343_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4551_ (.I(_0374_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4552_ (.A1(_3373_),
    .A2(_0372_),
    .A3(_0371_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4553_ (.A1(_0346_),
    .A2(_0371_),
    .A3(_0373_),
    .B1(_0375_),
    .B2(_0376_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4554_ (.A1(_3372_),
    .A2(_0178_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4555_ (.A1(_0377_),
    .A2(_0378_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4556_ (.A1(_0377_),
    .A2(_0378_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4557_ (.A1(_0345_),
    .A2(_0379_),
    .B(_0380_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4558_ (.A1(_0180_),
    .A2(_0241_),
    .A3(_3371_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4559_ (.A1(_0381_),
    .A2(_0382_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4560_ (.A1(_3297_),
    .A2(_2940_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4561_ (.A1(_3368_),
    .A2(_3174_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4562_ (.A1(_0306_),
    .A2(_0384_),
    .A3(_0385_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4563_ (.I(_0313_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4564_ (.A1(_0387_),
    .A2(_3075_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4565_ (.A1(_0385_),
    .A2(_0388_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4566_ (.A1(_0386_),
    .A2(_0389_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4567_ (.A1(_0387_),
    .A2(_0319_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4568_ (.I(\A[1][2] ),
    .Z(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4569_ (.A1(_0392_),
    .A2(_0971_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4570_ (.A1(_0314_),
    .A2(_2983_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4571_ (.I(_0392_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4572_ (.A1(_2983_),
    .A2(_0395_),
    .B1(_3072_),
    .B2(_3367_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4573_ (.A1(_0393_),
    .A2(_0394_),
    .B1(_0396_),
    .B2(_0384_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4574_ (.A1(_3310_),
    .A2(_0393_),
    .A3(_0308_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4575_ (.A1(_0397_),
    .A2(_0398_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4576_ (.A1(_0391_),
    .A2(_0399_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4577_ (.A1(_0390_),
    .A2(_0400_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4578_ (.A1(_0390_),
    .A2(_0400_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4579_ (.A1(_3015_),
    .A2(_0257_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4580_ (.A1(_0328_),
    .A2(_3098_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4581_ (.A1(_0282_),
    .A2(_3096_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4582_ (.A1(_0355_),
    .A2(_0404_),
    .A3(_0405_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4583_ (.I(_3101_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4584_ (.A1(_0351_),
    .A2(_0407_),
    .A3(_0350_),
    .A4(_3169_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4585_ (.A1(_0406_),
    .A2(_0408_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4586_ (.A1(_3043_),
    .A2(_3385_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4587_ (.I(_0152_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4588_ (.A1(_3101_),
    .A2(_0411_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4589_ (.A1(_0411_),
    .A2(_3043_),
    .B1(_0354_),
    .B2(_3039_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4590_ (.A1(_0410_),
    .A2(_0412_),
    .B1(_0413_),
    .B2(_0404_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4591_ (.A1(_3384_),
    .A2(_0410_),
    .A3(_0356_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4592_ (.A1(_0329_),
    .A2(_0414_),
    .A3(_0415_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4593_ (.A1(_0409_),
    .A2(_0416_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4594_ (.A1(_0409_),
    .A2(_0416_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4595_ (.A1(_0403_),
    .A2(_0417_),
    .B(_0418_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4596_ (.I(_3353_),
    .Z(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4597_ (.A1(_3007_),
    .A2(_0420_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4598_ (.A1(_0414_),
    .A2(_0415_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4599_ (.A1(_0414_),
    .A2(_0415_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4600_ (.A1(_0329_),
    .A2(_0422_),
    .B(_0423_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4601_ (.A1(_0330_),
    .A2(_0352_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4602_ (.A1(_0359_),
    .A2(_0360_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4603_ (.A1(_0425_),
    .A2(_0426_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4604_ (.A1(_0421_),
    .A2(_0424_),
    .A3(_0427_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4605_ (.A1(_0419_),
    .A2(_0428_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4606_ (.A1(_0419_),
    .A2(_0428_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4607_ (.A1(_0402_),
    .A2(_0429_),
    .B(_0430_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4608_ (.A1(_0321_),
    .A2(_0322_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4609_ (.A1(_0397_),
    .A2(_0398_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4610_ (.A1(_0341_),
    .A2(_0319_),
    .A3(_0399_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4611_ (.A1(_0433_),
    .A2(_0434_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4612_ (.A1(_0432_),
    .A2(_0435_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4613_ (.A1(_0424_),
    .A2(_0427_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4614_ (.A1(_0424_),
    .A2(_0427_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4615_ (.A1(_0421_),
    .A2(_0437_),
    .B(_0438_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4616_ (.A1(_0349_),
    .A2(_0365_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4617_ (.A1(_0436_),
    .A2(_0439_),
    .A3(_0440_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4618_ (.A1(_0431_),
    .A2(_0441_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4619_ (.A1(_0431_),
    .A2(_0441_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4620_ (.A1(_0401_),
    .A2(_0442_),
    .B(_0443_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4621_ (.A1(_0432_),
    .A2(_0435_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4622_ (.A1(_0315_),
    .A2(_0445_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4623_ (.A1(_0439_),
    .A2(_0440_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4624_ (.A1(_0439_),
    .A2(_0440_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4625_ (.A1(_0436_),
    .A2(_0447_),
    .B(_0448_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4626_ (.A1(_0347_),
    .A2(_0369_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4627_ (.A1(_0446_),
    .A2(_0449_),
    .A3(_0450_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4628_ (.A1(_0444_),
    .A2(_0451_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4629_ (.A1(_0316_),
    .A2(_0322_),
    .A3(_0435_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4630_ (.I(_0453_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4631_ (.A1(_0449_),
    .A2(_0450_),
    .Z(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4632_ (.A1(_0449_),
    .A2(_0450_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4633_ (.A1(_0446_),
    .A2(_0455_),
    .B(_0456_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4634_ (.A1(_0374_),
    .A2(_0376_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4635_ (.A1(_0454_),
    .A2(_0457_),
    .A3(_0458_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4636_ (.A1(_0419_),
    .A2(_0428_),
    .A3(_0402_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4637_ (.I(_0389_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4638_ (.A1(_0386_),
    .A2(_0461_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4639_ (.A1(_0406_),
    .A2(_0408_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4640_ (.A1(_3181_),
    .A2(_0190_),
    .A3(_0463_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4641_ (.A1(_0409_),
    .A2(_0416_),
    .A3(_0403_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4642_ (.A1(_0464_),
    .A2(_0465_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4643_ (.A1(_0464_),
    .A2(_0465_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4644_ (.A1(_0462_),
    .A2(_0466_),
    .B(_0467_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4645_ (.A1(_0460_),
    .A2(_0468_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4646_ (.I(_0469_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4647_ (.A1(_0464_),
    .A2(_0465_),
    .A3(_0462_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4648_ (.I(_3182_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4649_ (.I(_3369_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4650_ (.A1(_3181_),
    .A2(_0189_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4651_ (.A1(_0463_),
    .A2(_0474_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4652_ (.I(_0351_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4653_ (.A1(_0476_),
    .A2(_3169_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4654_ (.I(_0408_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4655_ (.A1(_0412_),
    .A2(_0477_),
    .B(_0478_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4656_ (.A1(_0472_),
    .A2(_0473_),
    .A3(_0475_),
    .A4(_0479_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4657_ (.A1(_0342_),
    .A2(_3174_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4658_ (.A1(_0394_),
    .A2(_0481_),
    .B(_0461_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4659_ (.A1(_3182_),
    .A2(_3369_),
    .A3(_0479_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4660_ (.A1(_0475_),
    .A2(_0483_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4661_ (.A1(_0482_),
    .A2(_0484_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4662_ (.A1(_0480_),
    .A2(_0485_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4663_ (.A1(_0471_),
    .A2(_0486_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4664_ (.A1(_3182_),
    .A2(_0473_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4665_ (.A1(_0479_),
    .A2(_0488_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4666_ (.I(_0476_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4667_ (.I(_0341_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4668_ (.A1(_0490_),
    .A2(_0491_),
    .A3(_0407_),
    .A4(_0472_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4669_ (.A1(_0489_),
    .A2(_0492_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4670_ (.A1(_0489_),
    .A2(_0492_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4671_ (.A1(_0388_),
    .A2(_0493_),
    .B(_0494_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4672_ (.A1(_0482_),
    .A2(_0484_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4673_ (.A1(_0495_),
    .A2(_0496_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4674_ (.A1(_0487_),
    .A2(_0497_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4675_ (.A1(_0470_),
    .A2(_0498_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4676_ (.A1(_0401_),
    .A2(_0431_),
    .A3(_0441_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4677_ (.A1(_0460_),
    .A2(_0468_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4678_ (.A1(_0480_),
    .A2(_0485_),
    .B(_0471_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4679_ (.A1(_0469_),
    .A2(_0502_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4680_ (.A1(_0501_),
    .A2(_0503_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4681_ (.A1(_0500_),
    .A2(_0504_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4682_ (.A1(_0499_),
    .A2(_0505_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4683_ (.A1(_0500_),
    .A2(_0503_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4684_ (.A1(_0444_),
    .A2(_0451_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4685_ (.A1(_0501_),
    .A2(_0500_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4686_ (.A1(_0508_),
    .A2(_0509_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4687_ (.A1(_0452_),
    .A2(_0459_),
    .B1(_0506_),
    .B2(_0507_),
    .C(_0510_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4688_ (.A1(_0508_),
    .A2(_0509_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4689_ (.A1(_0452_),
    .A2(_0512_),
    .B(_0459_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4690_ (.A1(_0511_),
    .A2(_0513_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4691_ (.A1(_0345_),
    .A2(_0379_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4692_ (.A1(_0457_),
    .A2(_0458_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4693_ (.A1(_0457_),
    .A2(_0458_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4694_ (.A1(_0454_),
    .A2(_0516_),
    .B(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4695_ (.A1(_0515_),
    .A2(_0518_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4696_ (.A1(_0383_),
    .A2(_0514_),
    .A3(_0519_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4697_ (.A1(_3371_),
    .A2(_0242_),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4698_ (.A1(_3371_),
    .A2(_0242_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4699_ (.A1(_0345_),
    .A2(_0379_),
    .B(_0382_),
    .C(_0380_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _4700_ (.A1(_0521_),
    .A2(_0381_),
    .A3(_0522_),
    .B1(_0523_),
    .B2(_0515_),
    .B3(_0518_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4701_ (.A1(_0520_),
    .A2(_0524_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4702_ (.A1(_0244_),
    .A2(_0301_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4703_ (.A1(_0304_),
    .A2(_0525_),
    .B(_0526_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4704_ (.A1(_0248_),
    .A2(_0299_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4705_ (.A1(_0246_),
    .A2(_0300_),
    .B(_0528_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4706_ (.I(_0257_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4707_ (.A1(_2909_),
    .A2(_0530_),
    .A3(_0254_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4708_ (.A1(_0250_),
    .A2(_0253_),
    .B(_0531_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4709_ (.A1(_0261_),
    .A2(_0297_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4710_ (.A1(_0259_),
    .A2(_0298_),
    .B(_0533_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4711_ (.A1(_1785_),
    .A2(_0420_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4712_ (.A1(_0289_),
    .A2(_0293_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4713_ (.A1(_0291_),
    .A2(_0536_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4714_ (.A1(_0285_),
    .A2(_0295_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4715_ (.A1(_0285_),
    .A2(_0295_),
    .Z(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4716_ (.A1(_0280_),
    .A2(_0538_),
    .B(_0539_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4717_ (.A1(_0537_),
    .A2(_0540_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4718_ (.A1(_0535_),
    .A2(_0541_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4719_ (.A1(_0263_),
    .A2(_0277_),
    .ZN(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4720_ (.A1(_0278_),
    .A2(_0296_),
    .B(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4721_ (.A1(_0208_),
    .A2(_0209_),
    .B1(_0288_),
    .B2(_0294_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4722_ (.I(_0220_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4723_ (.I(_0546_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4724_ (.I(_3383_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4725_ (.A1(_2930_),
    .A2(_3245_),
    .A3(_0547_),
    .A4(_0548_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4726_ (.A1(_0271_),
    .A2(_0274_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4727_ (.A1(_0549_),
    .A2(_0275_),
    .B(_0550_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4728_ (.A1(_0133_),
    .A2(_2942_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4729_ (.A1(_0286_),
    .A2(_0751_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4730_ (.A1(_0290_),
    .A2(_0553_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4731_ (.A1(_0552_),
    .A2(_0554_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4732_ (.A1(_0551_),
    .A2(_0555_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4733_ (.A1(_0545_),
    .A2(_0556_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4734_ (.A1(_0264_),
    .A2(_0268_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4735_ (.A1(_0269_),
    .A2(_0276_),
    .B(_0558_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4736_ (.A1(_0229_),
    .A2(_3033_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4737_ (.I(_0168_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4738_ (.I(_0561_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4739_ (.A1(_0562_),
    .A2(_3262_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4740_ (.A1(_0230_),
    .A2(_1235_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4741_ (.A1(_0265_),
    .A2(_0564_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4742_ (.A1(_0560_),
    .A2(_0563_),
    .B(_0565_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4743_ (.A1(_3393_),
    .A2(_2812_),
    .B1(_2813_),
    .B2(_0112_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4744_ (.A1(_0073_),
    .A2(_2969_),
    .A3(_2766_),
    .A4(_3380_),
    .Z(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4745_ (.A1(_0567_),
    .A2(_0568_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4746_ (.A1(_0265_),
    .A2(_0267_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4747_ (.A1(_0233_),
    .A2(_0560_),
    .B1(_0570_),
    .B2(_0266_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4748_ (.A1(_0569_),
    .A2(_0571_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4749_ (.A1(_0273_),
    .A2(_0572_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4750_ (.A1(_0566_),
    .A2(_0573_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4751_ (.A1(_0559_),
    .A2(_0574_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4752_ (.A1(_0557_),
    .A2(_0575_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4753_ (.A1(_0544_),
    .A2(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4754_ (.A1(_0542_),
    .A2(_0577_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4755_ (.A1(_0534_),
    .A2(_0578_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4756_ (.A1(_0532_),
    .A2(_0579_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4757_ (.A1(_0529_),
    .A2(_0580_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4758_ (.I(_0581_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4759_ (.A1(_0527_),
    .A2(_0582_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4760_ (.A1(_3295_),
    .A2(_0674_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4761_ (.I(_0584_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4762_ (.I(\B[2][6] ),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4763_ (.A1(_0586_),
    .A2(_1796_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4764_ (.I(\B[2][4] ),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4765_ (.A1(_1070_),
    .A2(_0588_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4766_ (.I(\B[2][5] ),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4767_ (.A1(_0590_),
    .A2(_0740_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4768_ (.A1(_0589_),
    .A2(_0591_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4769_ (.A1(_0587_),
    .A2(_0592_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4770_ (.I(\B[2][2] ),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4771_ (.A1(_1048_),
    .A2(_0594_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4772_ (.I(\B[2][1] ),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4773_ (.I(_0596_),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4774_ (.A1(_0597_),
    .A2(_0993_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4775_ (.I(\B[2][3] ),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4776_ (.I(_0599_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4777_ (.A1(_0600_),
    .A2(_0883_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4778_ (.A1(_1048_),
    .A2(_0596_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4779_ (.A1(_0594_),
    .A2(_0828_),
    .ZN(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4780_ (.A1(_0602_),
    .A2(_0603_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4781_ (.A1(_0595_),
    .A2(_0598_),
    .B1(_0601_),
    .B2(_0604_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4782_ (.A1(_1356_),
    .A2(_0596_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4783_ (.A1(_0600_),
    .A2(_0993_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4784_ (.A1(_0606_),
    .A2(_0595_),
    .A3(_0607_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4785_ (.A1(_0605_),
    .A2(_0608_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4786_ (.A1(_0605_),
    .A2(_0608_),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4787_ (.A1(_0593_),
    .A2(_0609_),
    .B(_0610_),
    .ZN(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4788_ (.I(\B[0][6] ),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4789_ (.I(_0612_),
    .Z(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4790_ (.A1(_0613_),
    .A2(_1323_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4791_ (.I(\B[2][0] ),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4792_ (.A1(_1378_),
    .A2(_0615_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4793_ (.A1(_0614_),
    .A2(_0616_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4794_ (.I(\B[0][4] ),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4795_ (.A1(_2201_),
    .A2(_0618_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4796_ (.I(\B[0][3] ),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4797_ (.A1(_2882_),
    .A2(_0620_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4798_ (.I(\B[0][5] ),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4799_ (.I(_0622_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4800_ (.A1(_0623_),
    .A2(_2931_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4801_ (.I(\B[0][3] ),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4802_ (.A1(_0625_),
    .A2(_2967_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4803_ (.I(\B[0][4] ),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4804_ (.I(_0627_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4805_ (.A1(_2810_),
    .A2(_0628_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4806_ (.A1(_0626_),
    .A2(_0629_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4807_ (.A1(_0619_),
    .A2(_0621_),
    .B1(_0624_),
    .B2(_0630_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4808_ (.A1(_2760_),
    .A2(\B[2][0] ),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4809_ (.I(\B[0][7] ),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4810_ (.A1(\B[0][6] ),
    .A2(_0633_),
    .A3(\A[2][0] ),
    .A4(_1180_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4811_ (.I(\B[0][6] ),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4812_ (.A1(_0633_),
    .A2(_1246_),
    .B1(_2814_),
    .B2(_0635_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4813_ (.A1(_0632_),
    .A2(_0634_),
    .A3(_0636_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4814_ (.A1(_0634_),
    .A2(_0636_),
    .B(_0632_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4815_ (.A1(_0637_),
    .A2(_0638_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4816_ (.A1(_0631_),
    .A2(_0639_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4817_ (.A1(_0631_),
    .A2(_0639_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4818_ (.A1(_0617_),
    .A2(_0640_),
    .B(_0641_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4819_ (.I(\B[2][6] ),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4820_ (.A1(_0643_),
    .A2(_2985_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4821_ (.A1(_0588_),
    .A2(_1532_),
    .ZN(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4822_ (.A1(_0590_),
    .A2(_1070_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4823_ (.A1(_0645_),
    .A2(_0646_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4824_ (.A1(_0644_),
    .A2(_0647_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4825_ (.I(\B[2][2] ),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4826_ (.A1(_1345_),
    .A2(_0649_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4827_ (.I(_0596_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4828_ (.I(_0594_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4829_ (.A1(_1367_),
    .A2(_0651_),
    .B1(_0652_),
    .B2(_2787_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4830_ (.A1(_0650_),
    .A2(_0602_),
    .B1(_0607_),
    .B2(_0653_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4831_ (.I(\B[2][1] ),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4832_ (.A1(_2790_),
    .A2(_0655_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4833_ (.A1(_2787_),
    .A2(_0599_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4834_ (.A1(_0650_),
    .A2(_0656_),
    .A3(_0657_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4835_ (.A1(_0654_),
    .A2(_0658_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4836_ (.A1(_0648_),
    .A2(_0659_),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4837_ (.A1(_0642_),
    .A2(_0660_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4838_ (.A1(_0642_),
    .A2(_0660_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4839_ (.A1(_0611_),
    .A2(_0661_),
    .B(_0662_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4840_ (.A1(_0590_),
    .A2(_0828_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4841_ (.A1(_0589_),
    .A2(_0664_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4842_ (.A1(_0644_),
    .A2(_0647_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4843_ (.A1(_0665_),
    .A2(_0666_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4844_ (.I(\B[2][7] ),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4845_ (.I(_0668_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4846_ (.I(_0669_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4847_ (.A1(_0663_),
    .A2(_0667_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4848_ (.A1(_0670_),
    .A2(_2910_),
    .A3(_0671_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4849_ (.A1(_0663_),
    .A2(_0667_),
    .B(_0672_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4850_ (.I(\B[2][7] ),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4851_ (.A1(_0675_),
    .A2(_2910_),
    .ZN(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4852_ (.A1(_0671_),
    .A2(_0676_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4853_ (.A1(_0642_),
    .A2(_0660_),
    .A3(_0611_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4854_ (.A1(_0617_),
    .A2(_0640_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4855_ (.A1(_0626_),
    .A2(_0629_),
    .A3(_0624_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4856_ (.I(\B[0][1] ),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4857_ (.I(_0681_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4858_ (.A1(_2157_),
    .A2(_0682_),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4859_ (.I(\B[0][0] ),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4860_ (.I(_0684_),
    .Z(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4861_ (.I(_0686_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4862_ (.A1(_0687_),
    .A2(_3271_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4863_ (.I(\B[0][2] ),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4864_ (.I(_0689_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4865_ (.A1(_0690_),
    .A2(_2806_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4866_ (.I(\B[0][1] ),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4867_ (.I(_0692_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4868_ (.I(_0693_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4869_ (.A1(_2452_),
    .A2(_0687_),
    .B1(_0694_),
    .B2(_2092_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4870_ (.A1(_0683_),
    .A2(_0688_),
    .B1(_0691_),
    .B2(_0695_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4871_ (.A1(_0689_),
    .A2(_2495_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4872_ (.I(_0684_),
    .Z(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4873_ (.A1(_3263_),
    .A2(_0699_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4874_ (.A1(_0683_),
    .A2(_0698_),
    .A3(_0700_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4875_ (.A1(_0697_),
    .A2(_0701_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4876_ (.A1(_0697_),
    .A2(_0701_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4877_ (.A1(_0680_),
    .A2(_0702_),
    .B(_0703_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4878_ (.A1(_0622_),
    .A2(_2882_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4879_ (.I(_0620_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4880_ (.A1(_0706_),
    .A2(_2092_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4881_ (.A1(_0619_),
    .A2(_0705_),
    .A3(_0708_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4882_ (.A1(_2704_),
    .A2(_0686_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4883_ (.A1(_2515_),
    .A2(_0681_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4884_ (.I(_0692_),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4885_ (.A1(_2525_),
    .A2(_0686_),
    .B1(_0712_),
    .B2(_2452_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4886_ (.A1(_0710_),
    .A2(_0711_),
    .B1(_0713_),
    .B2(_0698_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4887_ (.A1(_2146_),
    .A2(_0689_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4888_ (.I(\B[0][0] ),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4889_ (.A1(_2892_),
    .A2(_0716_),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _4890_ (.A1(_0711_),
    .A2(_0715_),
    .A3(_0717_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4891_ (.A1(_0714_),
    .A2(_0719_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4892_ (.A1(_0709_),
    .A2(_0720_),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4893_ (.A1(_0704_),
    .A2(_0721_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4894_ (.A1(_0704_),
    .A2(_0721_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4895_ (.A1(_0679_),
    .A2(_0722_),
    .B(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4896_ (.A1(_0632_),
    .A2(_0634_),
    .A3(_0636_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4897_ (.A1(_0634_),
    .A2(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4898_ (.A1(_0627_),
    .A2(_1949_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4899_ (.A1(_2967_),
    .A2(_0628_),
    .B1(_2430_),
    .B2(_0706_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _4900_ (.A1(_0626_),
    .A2(_0727_),
    .B1(_0728_),
    .B2(_0705_),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4901_ (.I(_0633_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4902_ (.A1(_0731_),
    .A2(_2354_),
    .B1(_2026_),
    .B2(_0612_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4903_ (.I(\B[0][6] ),
    .Z(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4904_ (.I(\B[0][7] ),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4905_ (.A1(_0733_),
    .A2(_0734_),
    .A3(_2814_),
    .A4(_2810_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4906_ (.A1(_0732_),
    .A2(_0735_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4907_ (.A1(_0730_),
    .A2(_0736_),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4908_ (.A1(_0726_),
    .A2(_0737_),
    .Z(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4909_ (.A1(_0714_),
    .A2(_0719_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4910_ (.A1(_0709_),
    .A2(_0720_),
    .B(_0739_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4911_ (.A1(_2892_),
    .A2(_0716_),
    .B1(_0682_),
    .B2(_2690_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4912_ (.A1(_2732_),
    .A2(_2821_),
    .A3(_0716_),
    .A4(_0682_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4913_ (.A1(_0715_),
    .A2(_0742_),
    .B(_0743_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4914_ (.A1(\A[2][7] ),
    .A2(_0681_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4915_ (.A1(_2515_),
    .A2(_0689_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4916_ (.A1(_0745_),
    .A2(_0746_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4917_ (.A1(_0744_),
    .A2(_0747_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4918_ (.A1(_2157_),
    .A2(\B[0][3] ),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4919_ (.A1(_0622_),
    .A2(_2201_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4920_ (.A1(_0727_),
    .A2(_0749_),
    .A3(_0750_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4921_ (.A1(_0748_),
    .A2(_0752_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4922_ (.A1(_0741_),
    .A2(_0753_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4923_ (.A1(_0738_),
    .A2(_0754_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4924_ (.A1(_0724_),
    .A2(_0755_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4925_ (.A1(_0724_),
    .A2(_0755_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4926_ (.A1(_0678_),
    .A2(_0756_),
    .B(_0757_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4927_ (.A1(_0648_),
    .A2(_0659_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4928_ (.A1(_0654_),
    .A2(_0658_),
    .B(_0759_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4929_ (.A1(_0730_),
    .A2(_0736_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4930_ (.A1(_0730_),
    .A2(_0736_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4931_ (.A1(_0726_),
    .A2(_0761_),
    .B(_0763_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4932_ (.A1(_0586_),
    .A2(_0883_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4933_ (.A1(_1444_),
    .A2(\B[2][4] ),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4934_ (.A1(_0664_),
    .A2(_0766_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4935_ (.A1(_0765_),
    .A2(_0767_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4936_ (.I(_0655_),
    .Z(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4937_ (.I(_0649_),
    .Z(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4938_ (.A1(_2937_),
    .A2(_0769_),
    .B1(_0770_),
    .B2(_1356_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4939_ (.A1(_2937_),
    .A2(_2785_),
    .A3(_0769_),
    .A4(_0770_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4940_ (.A1(_0771_),
    .A2(_0657_),
    .B(_0772_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4941_ (.A1(_2790_),
    .A2(_0649_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4942_ (.A1(_1499_),
    .A2(\B[2][3] ),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4943_ (.A1(_0775_),
    .A2(_0776_),
    .Z(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4944_ (.A1(_0774_),
    .A2(_0777_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4945_ (.A1(_0768_),
    .A2(_0778_),
    .Z(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4946_ (.A1(_0764_),
    .A2(_0779_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4947_ (.A1(_0760_),
    .A2(_0780_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4948_ (.A1(_0741_),
    .A2(_0753_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4949_ (.A1(_0738_),
    .A2(_0754_),
    .B(_0782_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4950_ (.A1(_2157_),
    .A2(\B[0][4] ),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4951_ (.A1(_0727_),
    .A2(_0749_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4952_ (.A1(_0708_),
    .A2(_0785_),
    .B1(_0786_),
    .B2(_0750_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4953_ (.A1(_0731_),
    .A2(_2026_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4954_ (.A1(_0733_),
    .A2(_2004_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4955_ (.A1(_0635_),
    .A2(_0734_),
    .A3(_2288_),
    .A4(_2267_),
    .Z(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4956_ (.A1(_0788_),
    .A2(_0789_),
    .B(_0790_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4957_ (.A1(_0787_),
    .A2(_0791_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4958_ (.A1(_0735_),
    .A2(_0792_),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4959_ (.A1(_0744_),
    .A2(_0747_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4960_ (.A1(_0748_),
    .A2(_0752_),
    .B(_0794_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4961_ (.A1(_0622_),
    .A2(_1949_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4962_ (.A1(_2690_),
    .A2(_0620_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _4963_ (.A1(_0785_),
    .A2(_0797_),
    .A3(_0798_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4964_ (.I(_0690_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4965_ (.A1(_3260_),
    .A2(_0800_),
    .A3(_0711_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4966_ (.A1(_0799_),
    .A2(_0801_),
    .Z(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4967_ (.A1(_0796_),
    .A2(_0802_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4968_ (.A1(_0793_),
    .A2(_0803_),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4969_ (.A1(_0783_),
    .A2(_0804_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4970_ (.A1(_0781_),
    .A2(_0805_),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4971_ (.A1(_0758_),
    .A2(_0807_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4972_ (.A1(_0758_),
    .A2(_0807_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4973_ (.A1(_0677_),
    .A2(_0808_),
    .B(_0809_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4974_ (.A1(_0760_),
    .A2(_0780_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4975_ (.A1(_0764_),
    .A2(_0779_),
    .B(_0811_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4976_ (.A1(_0664_),
    .A2(_0766_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4977_ (.A1(_0765_),
    .A2(_0767_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4978_ (.A1(_0813_),
    .A2(_0814_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4979_ (.A1(_0812_),
    .A2(_0815_),
    .Z(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4980_ (.A1(_0675_),
    .A2(_3225_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4981_ (.A1(_0816_),
    .A2(_0818_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4982_ (.A1(_0783_),
    .A2(_0804_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4983_ (.A1(_0781_),
    .A2(_0805_),
    .B(_0820_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4984_ (.A1(_0774_),
    .A2(_0777_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4985_ (.A1(_0768_),
    .A2(_0778_),
    .B(_0822_),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4986_ (.I(_0613_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4987_ (.A1(_0824_),
    .A2(_2933_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4988_ (.A1(_0787_),
    .A2(_0791_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4989_ (.A1(_0825_),
    .A2(_0788_),
    .A3(_0792_),
    .B(_0826_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4990_ (.I(_0599_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4991_ (.I(_0829_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4992_ (.A1(_2938_),
    .A2(_0830_),
    .A3(_0650_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4993_ (.A1(_0643_),
    .A2(_2943_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4994_ (.I(\B[2][5] ),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4995_ (.A1(_0833_),
    .A2(_2785_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4996_ (.A1(_0766_),
    .A2(_0834_),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4997_ (.I(_0833_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4998_ (.I(_0588_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4999_ (.A1(_0836_),
    .A2(_2949_),
    .B1(_0837_),
    .B2(_1367_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5000_ (.A1(_0835_),
    .A2(_0838_),
    .Z(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5001_ (.A1(_0832_),
    .A2(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5002_ (.A1(_0831_),
    .A2(_0841_),
    .Z(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5003_ (.A1(_0823_),
    .A2(_0827_),
    .A3(_0842_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5004_ (.A1(_0796_),
    .A2(_0802_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5005_ (.A1(_0793_),
    .A2(_0803_),
    .B(_0844_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5006_ (.A1(_0745_),
    .A2(_0746_),
    .B1(_0799_),
    .B2(_0801_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5007_ (.A1(_2525_),
    .A2(_0618_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5008_ (.I(\B[0][5] ),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5009_ (.A1(_0848_),
    .A2(_2452_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5010_ (.A1(_2893_),
    .A2(_0706_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5011_ (.A1(_0847_),
    .A2(_0849_),
    .A3(_0851_),
    .ZN(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5012_ (.A1(_0846_),
    .A2(_0852_),
    .ZN(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5013_ (.A1(_0785_),
    .A2(_0798_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5014_ (.A1(_0749_),
    .A2(_0847_),
    .B1(_0854_),
    .B2(_0797_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5015_ (.A1(_0734_),
    .A2(_2967_),
    .B1(_2092_),
    .B2(_0733_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5016_ (.A1(_0635_),
    .A2(_0633_),
    .A3(_2267_),
    .A4(_2660_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5017_ (.A1(_0856_),
    .A2(_0857_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5018_ (.A1(_0855_),
    .A2(_0858_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5019_ (.A1(_0790_),
    .A2(_0859_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5020_ (.A1(_0853_),
    .A2(_0860_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5021_ (.A1(_0845_),
    .A2(_0862_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5022_ (.A1(_0843_),
    .A2(_0863_),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5023_ (.A1(_0821_),
    .A2(_0864_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5024_ (.A1(_0819_),
    .A2(_0865_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5025_ (.A1(_0810_),
    .A2(_0866_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5026_ (.A1(_0673_),
    .A2(_0867_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5027_ (.A1(_0643_),
    .A2(_0718_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5028_ (.I(\B[2][4] ),
    .Z(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5029_ (.A1(_2984_),
    .A2(_0870_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5030_ (.A1(_0833_),
    .A2(_1576_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5031_ (.A1(_0871_),
    .A2(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5032_ (.A1(_0869_),
    .A2(_0874_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5033_ (.A1(_0651_),
    .A2(_0982_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5034_ (.A1(_0905_),
    .A2(_0829_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5035_ (.I(_0652_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5036_ (.A1(_0878_),
    .A2(_2922_),
    .B1(_2943_),
    .B2(_0597_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5037_ (.A1(_0603_),
    .A2(_0876_),
    .B1(_0877_),
    .B2(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5038_ (.A1(_0602_),
    .A2(_0603_),
    .A3(_0601_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5039_ (.A1(_0880_),
    .A2(_0881_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5040_ (.A1(_0880_),
    .A2(_0881_),
    .ZN(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5041_ (.A1(_0875_),
    .A2(_0882_),
    .B(_0884_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5042_ (.A1(_1180_),
    .A2(_0618_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5043_ (.A1(_0621_),
    .A2(_0886_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5044_ (.I(_0848_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5045_ (.A1(_0888_),
    .A2(_3008_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5046_ (.A1(_0621_),
    .A2(_0886_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5047_ (.A1(_0889_),
    .A2(_0890_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5048_ (.A1(_0614_),
    .A2(_0616_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5049_ (.A1(_0887_),
    .A2(_0891_),
    .B(_0892_),
    .C(_0617_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5050_ (.A1(_0605_),
    .A2(_0608_),
    .A3(_0593_),
    .Z(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5051_ (.A1(_0893_),
    .A2(_0895_),
    .Z(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5052_ (.A1(_0893_),
    .A2(_0895_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5053_ (.A1(_0885_),
    .A2(_0896_),
    .B(_0897_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5054_ (.A1(_0646_),
    .A2(_0871_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5055_ (.A1(_0587_),
    .A2(_0592_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5056_ (.A1(_0899_),
    .A2(_0900_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5057_ (.A1(_0898_),
    .A2(_0901_),
    .Z(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5058_ (.A1(_0898_),
    .A2(_0901_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5059_ (.A1(_0902_),
    .A2(_0903_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5060_ (.A1(_0675_),
    .A2(_1829_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5061_ (.A1(_0904_),
    .A2(_0906_),
    .B(_0902_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5062_ (.A1(_0904_),
    .A2(_0906_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5063_ (.A1(_0885_),
    .A2(_0896_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5064_ (.I(_0909_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5065_ (.A1(_0887_),
    .A2(_0891_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5066_ (.A1(_0617_),
    .A2(_0892_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5067_ (.A1(_0911_),
    .A2(_0912_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5068_ (.A1(_0889_),
    .A2(_0890_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5069_ (.A1(_0682_),
    .A2(_2081_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5070_ (.I(_0699_),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5071_ (.A1(_0917_),
    .A2(_3044_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5072_ (.A1(_0800_),
    .A2(_3108_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5073_ (.A1(_0694_),
    .A2(_3044_),
    .B1(_3271_),
    .B2(_0917_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5074_ (.A1(_0915_),
    .A2(_0918_),
    .B1(_0919_),
    .B2(_0920_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5075_ (.A1(_0710_),
    .A2(_0915_),
    .A3(_0691_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5076_ (.A1(_0921_),
    .A2(_0922_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5077_ (.A1(_0921_),
    .A2(_0922_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5078_ (.A1(_0914_),
    .A2(_0923_),
    .B(_0924_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5079_ (.A1(_0680_),
    .A2(_0702_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5080_ (.A1(_0925_),
    .A2(_0926_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5081_ (.A1(_0925_),
    .A2(_0926_),
    .Z(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5082_ (.A1(_0913_),
    .A2(_0928_),
    .B(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5083_ (.A1(_0704_),
    .A2(_0721_),
    .A3(_0679_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5084_ (.A1(_0930_),
    .A2(_0931_),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5085_ (.A1(_0913_),
    .A2(_0928_),
    .Z(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5086_ (.A1(_0929_),
    .A2(_0933_),
    .B(_0931_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5087_ (.A1(_0910_),
    .A2(_0932_),
    .B(_0934_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5088_ (.A1(_0678_),
    .A2(_0756_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5089_ (.A1(_0935_),
    .A2(_0936_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5090_ (.A1(_0935_),
    .A2(_0936_),
    .Z(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5091_ (.A1(_0908_),
    .A2(_0937_),
    .B(_0939_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5092_ (.A1(_0677_),
    .A2(_0808_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5093_ (.A1(_0940_),
    .A2(_0941_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5094_ (.A1(_0940_),
    .A2(_0941_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5095_ (.A1(_0907_),
    .A2(_0942_),
    .B(_0943_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5096_ (.A1(_0868_),
    .A2(_0944_),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5097_ (.I(_0770_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5098_ (.A1(_0946_),
    .A2(_0982_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5099_ (.I(_0597_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5100_ (.A1(_0948_),
    .A2(_2848_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5101_ (.I(_0600_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5102_ (.A1(_1796_),
    .A2(_0951_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5103_ (.I(_0946_),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5104_ (.A1(_0953_),
    .A2(_2848_),
    .B1(_2922_),
    .B2(_0948_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5105_ (.A1(_0947_),
    .A2(_0950_),
    .B1(_0952_),
    .B2(_0954_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5106_ (.A1(_0598_),
    .A2(_0947_),
    .A3(_0877_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5107_ (.A1(_0955_),
    .A2(_0956_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5108_ (.I(_0837_),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5109_ (.I(_0958_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5110_ (.A1(_2994_),
    .A2(_0959_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5111_ (.A1(_0873_),
    .A2(_0961_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5112_ (.I(_0836_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5113_ (.A1(_0963_),
    .A2(_2998_),
    .B1(_1818_),
    .B2(_0959_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5114_ (.A1(_0962_),
    .A2(_0964_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5115_ (.A1(_0955_),
    .A2(_0956_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5116_ (.A1(_0965_),
    .A2(_0966_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5117_ (.A1(_0957_),
    .A2(_0967_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5118_ (.I(_0615_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5119_ (.I(_0969_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5120_ (.I(_0625_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5121_ (.A1(_1323_),
    .A2(_0972_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5122_ (.A1(_0886_),
    .A2(_0973_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5123_ (.I(_0974_),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5124_ (.A1(_3005_),
    .A2(_0970_),
    .A3(_0975_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5125_ (.A1(_0875_),
    .A2(_0882_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5126_ (.A1(_0976_),
    .A2(_0977_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5127_ (.I(_3005_),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5128_ (.I(_0970_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5129_ (.A1(_0979_),
    .A2(_0980_),
    .A3(_0975_),
    .A4(_0977_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5130_ (.A1(_0968_),
    .A2(_0978_),
    .B(_0981_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5131_ (.A1(_0871_),
    .A2(_0873_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5132_ (.A1(_0869_),
    .A2(_0874_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5133_ (.A1(_0984_),
    .A2(_0985_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5134_ (.A1(_0983_),
    .A2(_0986_),
    .Z(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5135_ (.A1(_0983_),
    .A2(_0986_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5136_ (.A1(_0987_),
    .A2(_0988_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5137_ (.A1(_0675_),
    .A2(_3025_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5138_ (.A1(_0989_),
    .A2(_0990_),
    .B(_0987_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5139_ (.A1(_0910_),
    .A2(_0932_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5140_ (.A1(_0968_),
    .A2(_0978_),
    .Z(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5141_ (.A1(_3004_),
    .A2(_0970_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5142_ (.A1(_0975_),
    .A2(_0995_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5143_ (.I(_0625_),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5144_ (.I(_0997_),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5145_ (.I(_0628_),
    .Z(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5146_ (.I(_0999_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5147_ (.A1(_2933_),
    .A2(_0998_),
    .B1(_1000_),
    .B2(_3035_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5148_ (.I(_0693_),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5149_ (.A1(_1002_),
    .A2(_2004_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5150_ (.I(_0687_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5151_ (.A1(_1005_),
    .A2(_3246_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5152_ (.I(_0800_),
    .Z(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5153_ (.A1(_3106_),
    .A2(_1007_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5154_ (.I(_0712_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5155_ (.A1(_1009_),
    .A2(_3040_),
    .B1(_3247_),
    .B2(_1005_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5156_ (.A1(_1003_),
    .A2(_1006_),
    .B1(_1008_),
    .B2(_1010_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5157_ (.A1(_0688_),
    .A2(_1003_),
    .A3(_0919_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5158_ (.A1(_1011_),
    .A2(_1012_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5159_ (.A1(_1011_),
    .A2(_1012_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5160_ (.A1(_0975_),
    .A2(_1001_),
    .A3(_1013_),
    .B(_1014_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5161_ (.A1(_0914_),
    .A2(_0923_),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5162_ (.A1(_1016_),
    .A2(_1017_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5163_ (.A1(_1016_),
    .A2(_1017_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5164_ (.A1(_0996_),
    .A2(_1018_),
    .B(_1019_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5165_ (.A1(_0913_),
    .A2(_0928_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5166_ (.A1(_1020_),
    .A2(_1021_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5167_ (.A1(_1020_),
    .A2(_1021_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5168_ (.A1(_0994_),
    .A2(_1022_),
    .B(_1023_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5169_ (.A1(_0930_),
    .A2(_0931_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5170_ (.A1(_0909_),
    .A2(_1025_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5171_ (.A1(_0989_),
    .A2(_0990_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5172_ (.A1(_0909_),
    .A2(_1025_),
    .A3(_1024_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5173_ (.A1(_0992_),
    .A2(_1024_),
    .A3(_1027_),
    .B1(_1028_),
    .B2(_1029_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5174_ (.A1(_0908_),
    .A2(_0937_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5175_ (.A1(_1030_),
    .A2(_1031_),
    .Z(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5176_ (.A1(_1030_),
    .A2(_1031_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5177_ (.A1(_0991_),
    .A2(_1032_),
    .B(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5178_ (.A1(_0940_),
    .A2(_0941_),
    .A3(_0907_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5179_ (.A1(_1034_),
    .A2(_1035_),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5180_ (.A1(_0718_),
    .A2(_0951_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5181_ (.I(_0878_),
    .Z(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5182_ (.A1(_1807_),
    .A2(_1039_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5183_ (.A1(_0950_),
    .A2(_1038_),
    .A3(_1040_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5184_ (.I(_0651_),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5185_ (.I(_1042_),
    .Z(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5186_ (.A1(_2998_),
    .A2(_1043_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5187_ (.A1(_1040_),
    .A2(_1044_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5188_ (.A1(_1041_),
    .A2(_1045_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5189_ (.I(_0961_),
    .Z(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5190_ (.A1(_0652_),
    .A2(_2984_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5191_ (.A1(_1042_),
    .A2(_3081_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5192_ (.A1(_3081_),
    .A2(_0878_),
    .B1(_2848_),
    .B2(_1042_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5193_ (.A1(_1049_),
    .A2(_1050_),
    .B1(_1051_),
    .B2(_1038_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5194_ (.A1(_0876_),
    .A2(_1049_),
    .A3(_0952_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5195_ (.A1(_1052_),
    .A2(_1053_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5196_ (.A1(_1047_),
    .A2(_1054_),
    .Z(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5197_ (.A1(_1047_),
    .A2(_1054_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5198_ (.A1(_1046_),
    .A2(_1055_),
    .A3(_1056_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5199_ (.I(_1057_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5200_ (.A1(_1047_),
    .A2(_1046_),
    .A3(_1054_),
    .Z(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5201_ (.I(_1060_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5202_ (.I(_0969_),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5203_ (.A1(_1062_),
    .A2(_2923_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5204_ (.I(_1009_),
    .Z(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5205_ (.A1(_1064_),
    .A2(_2932_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5206_ (.A1(_3008_),
    .A2(_0800_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5207_ (.A1(_1006_),
    .A2(_1066_),
    .A3(_1065_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5208_ (.I(_0917_),
    .Z(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5209_ (.A1(_1068_),
    .A2(_3035_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5210_ (.A1(_1065_),
    .A2(_1067_),
    .A3(_1069_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5211_ (.A1(_1009_),
    .A2(_3108_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5212_ (.A1(_1005_),
    .A2(_3106_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5213_ (.A1(_1009_),
    .A2(_3106_),
    .B1(_3040_),
    .B2(_1005_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5214_ (.A1(_1072_),
    .A2(_1073_),
    .B1(_1074_),
    .B2(_1066_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5215_ (.A1(_0918_),
    .A2(_1072_),
    .A3(_1008_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5216_ (.A1(_0973_),
    .A2(_1075_),
    .A3(_1076_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5217_ (.A1(_1071_),
    .A2(_1077_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5218_ (.A1(_1071_),
    .A2(_1077_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5219_ (.A1(_1063_),
    .A2(_1078_),
    .B(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5220_ (.A1(_0970_),
    .A2(_3116_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5221_ (.A1(_1075_),
    .A2(_1076_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5222_ (.A1(_1075_),
    .A2(_1076_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5223_ (.A1(_0973_),
    .A2(_1083_),
    .B(_1084_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5224_ (.A1(_0974_),
    .A2(_1001_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5225_ (.A1(_1011_),
    .A2(_1012_),
    .Z(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5226_ (.A1(_1086_),
    .A2(_1087_),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5227_ (.A1(_1082_),
    .A2(_1085_),
    .A3(_1088_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5228_ (.A1(_1080_),
    .A2(_1089_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5229_ (.A1(_1080_),
    .A2(_1089_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5230_ (.A1(_1061_),
    .A2(_1090_),
    .B(_1091_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5231_ (.A1(_1052_),
    .A2(_1053_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5232_ (.A1(_1094_),
    .A2(_1055_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5233_ (.A1(_0965_),
    .A2(_0966_),
    .Z(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5234_ (.A1(_1095_),
    .A2(_1096_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5235_ (.A1(_1085_),
    .A2(_1088_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5236_ (.A1(_1085_),
    .A2(_1088_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5237_ (.A1(_1082_),
    .A2(_1098_),
    .B(_1099_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5238_ (.A1(_0996_),
    .A2(_1018_),
    .Z(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5239_ (.A1(_1097_),
    .A2(_1100_),
    .A3(_1101_),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5240_ (.A1(_1093_),
    .A2(_1102_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5241_ (.A1(_1093_),
    .A2(_1102_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5242_ (.A1(_1058_),
    .A2(_1104_),
    .B(_1105_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5243_ (.A1(_1095_),
    .A2(_1096_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5244_ (.A1(_0962_),
    .A2(_1107_),
    .Z(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5245_ (.A1(_1100_),
    .A2(_1101_),
    .Z(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5246_ (.A1(_1100_),
    .A2(_1101_),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5247_ (.A1(_1097_),
    .A2(_1109_),
    .B(_1110_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5248_ (.A1(_0994_),
    .A2(_1022_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5249_ (.A1(_1108_),
    .A2(_1111_),
    .A3(_1112_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5250_ (.A1(_1106_),
    .A2(_1113_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5251_ (.A1(_0873_),
    .A2(_1047_),
    .A3(_1107_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5252_ (.A1(_1111_),
    .A2(_1112_),
    .Z(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5253_ (.A1(_1111_),
    .A2(_1112_),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5254_ (.A1(_1108_),
    .A2(_1117_),
    .B(_1118_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5255_ (.A1(_1028_),
    .A2(_1029_),
    .Z(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5256_ (.A1(_1116_),
    .A2(_1119_),
    .A3(_1120_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5257_ (.A1(_1115_),
    .A2(_1121_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5258_ (.A1(_1057_),
    .A2(_1093_),
    .A3(_1102_),
    .Z(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5259_ (.A1(_1080_),
    .A2(_1089_),
    .A3(_1060_),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5260_ (.I(_1045_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5261_ (.A1(_1041_),
    .A2(_1126_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5262_ (.A1(_1065_),
    .A2(_1069_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5263_ (.A1(_1067_),
    .A2(_1128_),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5264_ (.A1(_1062_),
    .A2(_2849_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5265_ (.A1(_1129_),
    .A2(_1130_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5266_ (.A1(_1071_),
    .A2(_1077_),
    .A3(_1063_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5267_ (.A1(_1131_),
    .A2(_1132_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5268_ (.A1(_1131_),
    .A2(_1132_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5269_ (.A1(_1127_),
    .A2(_1133_),
    .B(_1134_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5270_ (.A1(_1124_),
    .A2(_1135_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5271_ (.A1(_1131_),
    .A2(_1132_),
    .A3(_1127_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5272_ (.A1(_1067_),
    .A2(_1128_),
    .A3(_1130_),
    .Z(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5273_ (.I(_1064_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5274_ (.A1(_3102_),
    .A2(_1140_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5275_ (.A1(_0980_),
    .A2(_1818_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5276_ (.A1(_1073_),
    .A2(_1141_),
    .B(_1142_),
    .C(_1128_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5277_ (.A1(_1139_),
    .A2(_1143_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5278_ (.A1(_3024_),
    .A2(_1039_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5279_ (.A1(_1050_),
    .A2(_1145_),
    .B(_1126_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5280_ (.A1(_1139_),
    .A2(_1143_),
    .Z(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5281_ (.A1(_1146_),
    .A2(_1148_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5282_ (.A1(_1144_),
    .A2(_1149_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5283_ (.A1(_1138_),
    .A2(_1150_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5284_ (.A1(_1137_),
    .A2(_1151_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5285_ (.A1(_1138_),
    .A2(_1150_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5286_ (.A1(_1073_),
    .A2(_1141_),
    .B(_1128_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5287_ (.A1(_1154_),
    .A2(_1142_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5288_ (.I(_1062_),
    .Z(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5289_ (.A1(_1156_),
    .A2(_3024_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5290_ (.A1(_1069_),
    .A2(_1157_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5291_ (.A1(_1155_),
    .A2(_1159_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5292_ (.A1(_1154_),
    .A2(_1142_),
    .A3(_1159_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5293_ (.A1(_1044_),
    .A2(_1161_),
    .Z(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5294_ (.A1(_1160_),
    .A2(_1162_),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5295_ (.A1(_1146_),
    .A2(_1148_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5296_ (.A1(_1163_),
    .A2(_1164_),
    .Z(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5297_ (.A1(_1153_),
    .A2(_1165_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5298_ (.A1(_1137_),
    .A2(_1166_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5299_ (.A1(_1124_),
    .A2(_1135_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5300_ (.A1(_1137_),
    .A2(_1151_),
    .B(_1168_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5301_ (.A1(_1123_),
    .A2(_1170_),
    .Z(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5302_ (.A1(_1167_),
    .A2(_1171_),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5303_ (.A1(_1123_),
    .A2(_1152_),
    .B(_1172_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5304_ (.A1(_1106_),
    .A2(_1113_),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5305_ (.A1(_1124_),
    .A2(_1135_),
    .A3(_1123_),
    .Z(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5306_ (.A1(_1174_),
    .A2(_1175_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5307_ (.A1(_1173_),
    .A2(_1176_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5308_ (.A1(_1174_),
    .A2(_1175_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5309_ (.A1(_1115_),
    .A2(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5310_ (.A1(_1119_),
    .A2(_1120_),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5311_ (.A1(_1116_),
    .A2(_1181_),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5312_ (.A1(_1122_),
    .A2(_1177_),
    .B1(_1179_),
    .B2(_1182_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5313_ (.A1(_0991_),
    .A2(_1032_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5314_ (.A1(_1119_),
    .A2(_1120_),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5315_ (.A1(_1116_),
    .A2(_1181_),
    .B(_1185_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5316_ (.A1(_1184_),
    .A2(_1186_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5317_ (.A1(_1036_),
    .A2(_1183_),
    .A3(_1187_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5318_ (.A1(_0907_),
    .A2(_0942_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5319_ (.A1(_0907_),
    .A2(_0942_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5320_ (.A1(_0991_),
    .A2(_1032_),
    .B(_1035_),
    .C(_1033_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _5321_ (.A1(_1189_),
    .A2(_1034_),
    .A3(_1190_),
    .B1(_1192_),
    .B2(_1184_),
    .B3(_1186_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5322_ (.A1(_0868_),
    .A2(_0944_),
    .Z(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5323_ (.A1(_1188_),
    .A2(_1193_),
    .B(_1194_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5324_ (.A1(_0945_),
    .A2(_1195_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5325_ (.A1(_0810_),
    .A2(_0866_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5326_ (.A1(_0673_),
    .A2(_0867_),
    .B(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5327_ (.I(_0668_),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5328_ (.I(_1199_),
    .Z(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5329_ (.A1(_1200_),
    .A2(_3225_),
    .A3(_0816_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5330_ (.A1(_0812_),
    .A2(_0815_),
    .B(_1201_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5331_ (.I(_1203_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5332_ (.A1(_0821_),
    .A2(_0864_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5333_ (.A1(_0819_),
    .A2(_0865_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5334_ (.A1(_1205_),
    .A2(_1206_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5335_ (.I(_3116_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5336_ (.A1(_1199_),
    .A2(_1208_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5337_ (.A1(_0832_),
    .A2(_0840_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5338_ (.A1(_0835_),
    .A2(_1210_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5339_ (.A1(_0827_),
    .A2(_0842_),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5340_ (.A1(_0827_),
    .A2(_0842_),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5341_ (.A1(_0823_),
    .A2(_1212_),
    .B(_1214_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5342_ (.A1(_1211_),
    .A2(_1215_),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5343_ (.A1(_1209_),
    .A2(_1216_),
    .Z(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5344_ (.A1(_0845_),
    .A2(_0862_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5345_ (.A1(_0843_),
    .A2(_0863_),
    .B(_1218_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5346_ (.A1(_0775_),
    .A2(_0776_),
    .B1(_0831_),
    .B2(_0841_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5347_ (.I(_0734_),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5348_ (.I(_1221_),
    .Z(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5349_ (.I(_1222_),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5350_ (.A1(_0824_),
    .A2(_1223_),
    .A3(_3246_),
    .A4(_3247_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5351_ (.A1(_0855_),
    .A2(_0858_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5352_ (.A1(_1225_),
    .A2(_0859_),
    .B(_1226_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5353_ (.I(_0586_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5354_ (.I(_1228_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5355_ (.A1(_1229_),
    .A2(_3004_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5356_ (.A1(_2938_),
    .A2(_0958_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5357_ (.A1(_0834_),
    .A2(_1231_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5358_ (.A1(_1230_),
    .A2(_1232_),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5359_ (.A1(_1227_),
    .A2(_1233_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5360_ (.A1(_1220_),
    .A2(_1234_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5361_ (.A1(_0846_),
    .A2(_0852_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5362_ (.A1(_0853_),
    .A2(_0860_),
    .B(_1237_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5363_ (.I(_2893_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5364_ (.A1(_1239_),
    .A2(_0999_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5365_ (.I(_0888_),
    .Z(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5366_ (.A1(_1241_),
    .A2(_3264_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5367_ (.A1(_0888_),
    .A2(_3260_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5368_ (.A1(_0847_),
    .A2(_1243_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5369_ (.A1(_1240_),
    .A2(_1242_),
    .B(_1244_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5370_ (.I(_0612_),
    .Z(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5371_ (.I(_0731_),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5372_ (.A1(_1247_),
    .A2(_3270_),
    .B1(_3272_),
    .B2(_1248_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5373_ (.I(_0733_),
    .Z(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5374_ (.A1(_1250_),
    .A2(_1248_),
    .A3(_3270_),
    .A4(_3272_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5375_ (.A1(_1249_),
    .A2(_1251_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5376_ (.A1(_0847_),
    .A2(_0851_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5377_ (.A1(_0798_),
    .A2(_1240_),
    .B1(_1253_),
    .B2(_0849_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5378_ (.A1(_1252_),
    .A2(_1254_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5379_ (.A1(_0857_),
    .A2(_1255_),
    .Z(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5380_ (.A1(_1245_),
    .A2(_1256_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5381_ (.A1(_1238_),
    .A2(_1258_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5382_ (.A1(_1236_),
    .A2(_1259_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5383_ (.A1(_1219_),
    .A2(_1260_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5384_ (.A1(_1217_),
    .A2(_1261_),
    .Z(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5385_ (.A1(_1204_),
    .A2(_1207_),
    .A3(_1262_),
    .Z(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5386_ (.A1(_1198_),
    .A2(_1263_),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5387_ (.A1(_1196_),
    .A2(_1264_),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5388_ (.A1(_3296_),
    .A2(_0583_),
    .B1(_0585_),
    .B2(_1265_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5389_ (.I(net2),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5390_ (.I(_1267_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5391_ (.I(_1269_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5392_ (.I(_3289_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5393_ (.A1(_3295_),
    .A2(_1271_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5394_ (.I(_1272_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5395_ (.I(_1273_),
    .Z(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5396_ (.A1(_1247_),
    .A2(_3328_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5397_ (.A1(_3334_),
    .A2(_0615_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5398_ (.A1(_1275_),
    .A2(_1276_),
    .Z(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5399_ (.I(_0627_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5400_ (.A1(_0149_),
    .A2(_1278_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5401_ (.A1(\A[0][2] ),
    .A2(_0620_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5402_ (.A1(_0161_),
    .A2(_0625_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5403_ (.A1(_3399_),
    .A2(_0618_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5404_ (.A1(_1282_),
    .A2(_1283_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5405_ (.A1(_0623_),
    .A2(_0065_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5406_ (.A1(_1280_),
    .A2(_1281_),
    .B1(_1284_),
    .B2(_1285_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5407_ (.A1(_0286_),
    .A2(_0615_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5408_ (.A1(_0635_),
    .A2(_3325_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5409_ (.A1(_0731_),
    .A2(_0327_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5410_ (.A1(_1287_),
    .A2(_1288_),
    .A3(_1289_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5411_ (.A1(_1286_),
    .A2(_1291_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5412_ (.A1(_1277_),
    .A2(_1292_),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5413_ (.A1(\A[0][5] ),
    .A2(_0681_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5414_ (.A1(_0686_),
    .A2(_0069_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5415_ (.I(\B[0][2] ),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5416_ (.A1(_1296_),
    .A2(_3390_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5417_ (.A1(_0073_),
    .A2(_0699_),
    .B1(_0712_),
    .B2(_3380_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5418_ (.A1(_1294_),
    .A2(_1295_),
    .B1(_1297_),
    .B2(_1298_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5419_ (.A1(\A[0][6] ),
    .A2(\B[0][0] ),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5420_ (.A1(_1296_),
    .A2(_0111_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5421_ (.A1(_1294_),
    .A2(_1300_),
    .A3(_1302_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5422_ (.A1(_1299_),
    .A2(_1303_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5423_ (.A1(_1282_),
    .A2(_1283_),
    .A3(_1285_),
    .Z(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5424_ (.A1(_1299_),
    .A2(_1303_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5425_ (.A1(_1304_),
    .A2(_1305_),
    .B(_1306_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5426_ (.A1(_0072_),
    .A2(_0684_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5427_ (.A1(_0102_),
    .A2(_0692_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5428_ (.I(_0716_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5429_ (.I(_3392_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5430_ (.A1(_0080_),
    .A2(_1310_),
    .B1(_1002_),
    .B2(_1311_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5431_ (.A1(_1308_),
    .A2(_1309_),
    .B1(_1313_),
    .B2(_1302_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5432_ (.A1(_0164_),
    .A2(_0684_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5433_ (.A1(_0073_),
    .A2(_1296_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5434_ (.A1(_1309_),
    .A2(_1315_),
    .A3(_1316_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5435_ (.A1(_1314_),
    .A2(_1317_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5436_ (.A1(_0848_),
    .A2(_0220_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5437_ (.A1(_0997_),
    .A2(_3387_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5438_ (.A1(_1280_),
    .A2(_1319_),
    .A3(_1320_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5439_ (.A1(_1318_),
    .A2(_1321_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5440_ (.A1(_1307_),
    .A2(_1322_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5441_ (.A1(_1293_),
    .A2(_1324_),
    .Z(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5442_ (.A1(\A[0][1] ),
    .A2(_0627_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5443_ (.A1(_1281_),
    .A2(_1326_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5444_ (.A1(_0623_),
    .A2(_0327_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5445_ (.A1(_1281_),
    .A2(_1326_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5446_ (.A1(_1328_),
    .A2(_1329_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5447_ (.A1(_1327_),
    .A2(_1330_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5448_ (.A1(_1275_),
    .A2(_1276_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5449_ (.A1(_1277_),
    .A2(_1332_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5450_ (.A1(_1331_),
    .A2(_1333_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5451_ (.A1(_1328_),
    .A2(_1329_),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5452_ (.A1(_0692_),
    .A2(_3379_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5453_ (.A1(_1310_),
    .A2(_0088_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5454_ (.A1(_3323_),
    .A2(_0690_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5455_ (.A1(_1002_),
    .A2(_0161_),
    .B1(_0112_),
    .B2(_0699_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5456_ (.A1(_1337_),
    .A2(_1338_),
    .B1(_1339_),
    .B2(_1340_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5457_ (.A1(_1308_),
    .A2(_1337_),
    .A3(_1297_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5458_ (.A1(_1341_),
    .A2(_1342_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5459_ (.A1(_1341_),
    .A2(_1342_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5460_ (.A1(_1336_),
    .A2(_1343_),
    .B(_1344_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5461_ (.A1(_1304_),
    .A2(_1305_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5462_ (.A1(_1346_),
    .A2(_1347_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5463_ (.A1(_1346_),
    .A2(_1347_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5464_ (.A1(_1335_),
    .A2(_1348_),
    .B(_1349_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5465_ (.A1(_1293_),
    .A2(_1324_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5466_ (.A1(_0586_),
    .A2(\A[1][0] ),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5467_ (.A1(\A[1][2] ),
    .A2(_0588_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5468_ (.A1(_0590_),
    .A2(\A[1][1] ),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5469_ (.A1(_1353_),
    .A2(_1354_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5470_ (.A1(_1352_),
    .A2(_1355_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5471_ (.A1(_0649_),
    .A2(\A[1][4] ),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5472_ (.A1(_0651_),
    .A2(_3317_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5473_ (.A1(_0652_),
    .A2(_3308_),
    .B1(_3305_),
    .B2(_0769_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5474_ (.A1(_3299_),
    .A2(_0600_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5475_ (.A1(_1358_),
    .A2(_1359_),
    .B1(_1360_),
    .B2(_1361_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5476_ (.A1(\A[1][5] ),
    .A2(_0655_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5477_ (.A1(\A[1][3] ),
    .A2(_0599_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5478_ (.A1(_1363_),
    .A2(_1358_),
    .A3(_1364_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5479_ (.A1(_1362_),
    .A2(_1365_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5480_ (.A1(_1362_),
    .A2(_1365_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5481_ (.A1(_1357_),
    .A2(_1366_),
    .B(_1368_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5482_ (.A1(_1327_),
    .A2(_1330_),
    .B(_1332_),
    .C(_1277_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5483_ (.A1(_3345_),
    .A2(_0770_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5484_ (.A1(_0597_),
    .A2(_0128_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5485_ (.A1(_1363_),
    .A2(_1358_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5486_ (.A1(_1371_),
    .A2(_1372_),
    .B1(_1373_),
    .B2(_1364_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5487_ (.A1(_3333_),
    .A2(_0769_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5488_ (.A1(_0829_),
    .A2(_0128_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5489_ (.A1(_1375_),
    .A2(_1371_),
    .A3(_1376_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5490_ (.A1(_0643_),
    .A2(_0307_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5491_ (.I(_0833_),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5492_ (.A1(_1380_),
    .A2(_3299_),
    .A3(_3317_),
    .A4(_0870_),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5493_ (.A1(_1380_),
    .A2(_0392_),
    .B1(_0255_),
    .B2(_0837_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5494_ (.A1(_1381_),
    .A2(_1382_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5495_ (.A1(_1379_),
    .A2(_1383_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5496_ (.A1(_1374_),
    .A2(_1377_),
    .A3(_1384_),
    .Z(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5497_ (.A1(_1370_),
    .A2(_1385_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5498_ (.A1(_1369_),
    .A2(_1386_),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5499_ (.I(_1387_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5500_ (.A1(_1293_),
    .A2(_1324_),
    .Z(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5501_ (.A1(_1350_),
    .A2(_1390_),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5502_ (.A1(_1325_),
    .A2(_1350_),
    .A3(_1351_),
    .B1(_1388_),
    .B2(_1391_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5503_ (.A1(_1286_),
    .A2(_1291_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5504_ (.A1(_1277_),
    .A2(_1292_),
    .B(_1393_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5505_ (.A1(_1228_),
    .A2(_3311_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5506_ (.A1(_1380_),
    .A2(_0255_),
    .A3(_0128_),
    .A4(_0870_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5507_ (.A1(_0836_),
    .A2(_3309_),
    .B1(_3313_),
    .B2(_0837_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5508_ (.A1(_1396_),
    .A2(_1397_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5509_ (.A1(_1395_),
    .A2(_1398_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5510_ (.A1(_3350_),
    .A2(_0594_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5511_ (.A1(_1375_),
    .A2(_1371_),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5512_ (.A1(_1401_),
    .A2(_1363_),
    .B1(_1402_),
    .B2(_1376_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5513_ (.A1(_0136_),
    .A2(_0655_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5514_ (.A1(_1401_),
    .A2(_1404_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5515_ (.A1(_3346_),
    .A2(_0829_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5516_ (.A1(_1405_),
    .A2(_1406_),
    .Z(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5517_ (.A1(_1403_),
    .A2(_1407_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5518_ (.A1(_1399_),
    .A2(_1408_),
    .Z(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5519_ (.A1(_1374_),
    .A2(_1377_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5520_ (.A1(_1374_),
    .A2(_1377_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5521_ (.A1(_1384_),
    .A2(_1410_),
    .B(_1412_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5522_ (.A1(_1394_),
    .A2(_1409_),
    .A3(_1413_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5523_ (.A1(_1307_),
    .A2(_1322_),
    .Z(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5524_ (.A1(_1293_),
    .A2(_1324_),
    .B(_1415_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5525_ (.A1(_1314_),
    .A2(_1317_),
    .ZN(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5526_ (.A1(_1318_),
    .A2(_1321_),
    .B(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5527_ (.A1(_0229_),
    .A2(_1310_),
    .B1(_0712_),
    .B2(_0168_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5528_ (.A1(_0229_),
    .A2(_0168_),
    .A3(_1310_),
    .A4(_1002_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5529_ (.A1(_1419_),
    .A2(_1316_),
    .B(_1420_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5530_ (.A1(_0164_),
    .A2(_0693_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5531_ (.A1(_0079_),
    .A2(_1296_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5532_ (.A1(_1423_),
    .A2(_1424_),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5533_ (.A1(_1421_),
    .A2(_1425_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5534_ (.A1(_0112_),
    .A2(_0628_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5535_ (.A1(_0848_),
    .A2(_0088_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5536_ (.A1(_1311_),
    .A2(_0997_),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5537_ (.A1(_1427_),
    .A2(_1428_),
    .A3(_1429_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5538_ (.A1(_1426_),
    .A2(_1430_),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5539_ (.A1(_1418_),
    .A2(_1431_),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5540_ (.A1(_1248_),
    .A2(_0281_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5541_ (.A1(_1288_),
    .A2(_1289_),
    .Z(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5542_ (.A1(_1275_),
    .A2(_1434_),
    .B1(_1435_),
    .B2(_1287_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5543_ (.I(_0070_),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5544_ (.A1(_0972_),
    .A2(_1437_),
    .B1(_0999_),
    .B2(_0357_),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5545_ (.A1(_1282_),
    .A2(_1427_),
    .B1(_1438_),
    .B2(_1319_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5546_ (.A1(_1247_),
    .A2(_0546_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5547_ (.A1(_1250_),
    .A2(_1221_),
    .A3(_0152_),
    .A4(_0546_),
    .Z(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5548_ (.A1(_1434_),
    .A2(_1440_),
    .B(_1441_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5549_ (.A1(_1439_),
    .A2(_1442_),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5550_ (.A1(_1436_),
    .A2(_1443_),
    .Z(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5551_ (.A1(_1432_),
    .A2(_1445_),
    .Z(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5552_ (.A1(_1416_),
    .A2(_1446_),
    .Z(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5553_ (.A1(_1414_),
    .A2(_1447_),
    .Z(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5554_ (.A1(_1392_),
    .A2(_1448_),
    .Z(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5555_ (.A1(_1370_),
    .A2(_1385_),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5556_ (.A1(_1369_),
    .A2(_1386_),
    .B(_1450_),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5557_ (.A1(_1379_),
    .A2(_1383_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5558_ (.A1(_1381_),
    .A2(_1452_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5559_ (.A1(_1451_),
    .A2(_1453_),
    .Z(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5560_ (.A1(_1451_),
    .A2(_1453_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5561_ (.A1(_1454_),
    .A2(_1456_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5562_ (.A1(_0668_),
    .A2(_0473_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5563_ (.A1(_1457_),
    .A2(_1458_),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5564_ (.A1(_1392_),
    .A2(_1448_),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5565_ (.A1(_1459_),
    .A2(_1460_),
    .Z(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5566_ (.A1(_1394_),
    .A2(_1409_),
    .Z(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5567_ (.A1(_1394_),
    .A2(_1409_),
    .Z(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5568_ (.A1(_1413_),
    .A2(_1462_),
    .B(_1463_),
    .ZN(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5569_ (.A1(_1395_),
    .A2(_1398_),
    .ZN(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5570_ (.A1(_1396_),
    .A2(_1465_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5571_ (.A1(_1464_),
    .A2(_1467_),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5572_ (.A1(_0669_),
    .A2(_0191_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5573_ (.A1(_1468_),
    .A2(_1469_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5574_ (.A1(_1415_),
    .A2(_1325_),
    .B(_1446_),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5575_ (.A1(_1414_),
    .A2(_1447_),
    .B(_1471_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5576_ (.A1(_1418_),
    .A2(_1431_),
    .Z(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5577_ (.A1(_1432_),
    .A2(_1445_),
    .B(_1473_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5578_ (.A1(_1421_),
    .A2(_1425_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5579_ (.A1(_1426_),
    .A2(_1430_),
    .B(_1475_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5580_ (.A1(_1311_),
    .A2(_1278_),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5581_ (.A1(_0623_),
    .A2(_0070_),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5582_ (.A1(_0561_),
    .A2(_0972_),
    .ZN(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5583_ (.A1(_1478_),
    .A2(_1479_),
    .A3(_1480_),
    .Z(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5584_ (.I(_0230_),
    .Z(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5585_ (.A1(_1482_),
    .A2(_1007_),
    .A3(_1309_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5586_ (.A1(_1481_),
    .A2(_1483_),
    .Z(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5587_ (.A1(_1476_),
    .A2(_1484_),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5588_ (.I(_0075_),
    .Z(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5589_ (.A1(_1486_),
    .A2(_0998_),
    .B1(_1437_),
    .B2(_0999_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5590_ (.A1(_1320_),
    .A2(_1478_),
    .B1(_1487_),
    .B2(_1428_),
    .ZN(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5591_ (.A1(_0613_),
    .A2(_1222_),
    .A3(_0354_),
    .A4(_0357_),
    .Z(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5592_ (.A1(_1222_),
    .A2(_0547_),
    .B1(_0548_),
    .B2(_0613_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5593_ (.A1(_1490_),
    .A2(_1491_),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5594_ (.A1(_1489_),
    .A2(_1492_),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5595_ (.A1(_1441_),
    .A2(_1493_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5596_ (.A1(_1485_),
    .A2(_1494_),
    .Z(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5597_ (.A1(_1474_),
    .A2(_1495_),
    .Z(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5598_ (.A1(_1403_),
    .A2(_1407_),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5599_ (.A1(_1399_),
    .A2(_1408_),
    .B(_1497_),
    .ZN(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5600_ (.A1(_1439_),
    .A2(_1442_),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5601_ (.A1(_1436_),
    .A2(_1443_),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5602_ (.A1(_1500_),
    .A2(_1501_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5603_ (.A1(_1228_),
    .A2(_0256_),
    .ZN(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5604_ (.A1(_1380_),
    .A2(_3313_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5605_ (.A1(_3346_),
    .A2(_0870_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5606_ (.A1(_1504_),
    .A2(_1505_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5607_ (.A1(_1503_),
    .A2(_1506_),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5608_ (.A1(_0286_),
    .A2(_0878_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5609_ (.A1(_1375_),
    .A2(_1508_),
    .B1(_1405_),
    .B2(_1406_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5610_ (.A1(_3351_),
    .A2(_0951_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5611_ (.A1(_1508_),
    .A2(_1511_),
    .Z(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5612_ (.A1(_1509_),
    .A2(_1512_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5613_ (.A1(_1507_),
    .A2(_1513_),
    .Z(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5614_ (.A1(_1502_),
    .A2(_1514_),
    .Z(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5615_ (.A1(_1498_),
    .A2(_1515_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5616_ (.A1(_1496_),
    .A2(_1516_),
    .Z(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5617_ (.A1(_1472_),
    .A2(_1517_),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5618_ (.A1(_1470_),
    .A2(_1518_),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5619_ (.A1(_1449_),
    .A2(_1461_),
    .B(_1519_),
    .ZN(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5620_ (.A1(_1457_),
    .A2(_1458_),
    .B(_1454_),
    .ZN(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5621_ (.A1(_1459_),
    .A2(_1460_),
    .B(_1449_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5622_ (.A1(_1523_),
    .A2(_1519_),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5623_ (.A1(_1522_),
    .A2(_1524_),
    .ZN(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5624_ (.I(_1200_),
    .Z(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5625_ (.A1(_1526_),
    .A2(_0191_),
    .A3(_1468_),
    .ZN(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5626_ (.A1(_1464_),
    .A2(_1467_),
    .B(_1527_),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5627_ (.A1(_1472_),
    .A2(_1517_),
    .Z(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5628_ (.A1(_1470_),
    .A2(_1518_),
    .B(_1529_),
    .ZN(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5629_ (.A1(_1432_),
    .A2(_1445_),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5630_ (.A1(_1473_),
    .A2(_1531_),
    .B(_1495_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5631_ (.A1(_1496_),
    .A2(_1516_),
    .B(_1533_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5632_ (.A1(_1476_),
    .A2(_1484_),
    .ZN(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5633_ (.A1(_1485_),
    .A2(_1494_),
    .B(_1535_),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5634_ (.A1(_1423_),
    .A2(_1424_),
    .B1(_1481_),
    .B2(_1483_),
    .ZN(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5635_ (.A1(_1241_),
    .A2(_1486_),
    .ZN(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5636_ (.A1(_0080_),
    .A2(_1278_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5637_ (.A1(_0230_),
    .A2(_0706_),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5638_ (.A1(_1539_),
    .A2(_1540_),
    .ZN(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5639_ (.A1(_1538_),
    .A2(_1541_),
    .Z(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5640_ (.A1(_1537_),
    .A2(_1542_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5641_ (.A1(_0824_),
    .A2(_1223_),
    .A3(_0547_),
    .A4(_0548_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5642_ (.A1(_1248_),
    .A2(_0357_),
    .ZN(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5643_ (.A1(_0561_),
    .A2(_0997_),
    .B1(_1278_),
    .B2(_1311_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5644_ (.A1(_1429_),
    .A2(_1539_),
    .B1(_1547_),
    .B2(_1479_),
    .ZN(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5645_ (.A1(_0612_),
    .A2(_3387_),
    .ZN(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5646_ (.A1(_1546_),
    .A2(_1548_),
    .A3(_1549_),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5647_ (.A1(_1545_),
    .A2(_1550_),
    .Z(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5648_ (.A1(_1544_),
    .A2(_1551_),
    .Z(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5649_ (.A1(_1536_),
    .A2(_1552_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5650_ (.A1(_1509_),
    .A2(_1512_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5651_ (.A1(_1507_),
    .A2(_1513_),
    .B(_1555_),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5652_ (.A1(_1489_),
    .A2(_1492_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5653_ (.A1(_1441_),
    .A2(_1493_),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5654_ (.A1(_1557_),
    .A2(_1558_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5655_ (.A1(_0287_),
    .A2(_0830_),
    .A3(_1401_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5656_ (.A1(_1228_),
    .A2(_3353_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5657_ (.A1(_0836_),
    .A2(_3334_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5658_ (.A1(_1505_),
    .A2(_1562_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5659_ (.I(_3334_),
    .Z(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5660_ (.A1(_0963_),
    .A2(_0133_),
    .B1(_0958_),
    .B2(_1564_),
    .ZN(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5661_ (.A1(_1563_),
    .A2(_1566_),
    .Z(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5662_ (.A1(_1561_),
    .A2(_1567_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5663_ (.A1(_1560_),
    .A2(_1568_),
    .Z(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5664_ (.A1(_1556_),
    .A2(_1559_),
    .A3(_1569_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5665_ (.A1(_1553_),
    .A2(_1570_),
    .Z(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5666_ (.A1(_1502_),
    .A2(_1514_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5667_ (.A1(_1498_),
    .A2(_1515_),
    .B(_1572_),
    .ZN(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5668_ (.A1(_1504_),
    .A2(_1505_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5669_ (.A1(_1503_),
    .A2(_1506_),
    .ZN(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5670_ (.A1(_1574_),
    .A2(_1575_),
    .ZN(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5671_ (.A1(_1573_),
    .A2(_1577_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5672_ (.A1(_1199_),
    .A2(_0530_),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5673_ (.A1(_1578_),
    .A2(_1579_),
    .Z(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5674_ (.A1(_1534_),
    .A2(_1571_),
    .A3(_1580_),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5675_ (.A1(_1530_),
    .A2(_1581_),
    .ZN(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5676_ (.A1(_1528_),
    .A2(_1582_),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5677_ (.A1(_1520_),
    .A2(_1525_),
    .B(_1583_),
    .ZN(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5678_ (.A1(_1520_),
    .A2(_1525_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5679_ (.A1(_1583_),
    .A2(_1585_),
    .ZN(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5680_ (.A1(_0946_),
    .A2(_0255_),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5681_ (.A1(_0948_),
    .A2(_0395_),
    .ZN(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5682_ (.A1(_0395_),
    .A2(_0953_),
    .B1(_0256_),
    .B2(_1042_),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5683_ (.A1(_0307_),
    .A2(_0951_),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5684_ (.A1(_1588_),
    .A2(_1589_),
    .B1(_1590_),
    .B2(_1591_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5685_ (.A1(_1372_),
    .A2(_1588_),
    .A3(_1361_),
    .ZN(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5686_ (.A1(_1592_),
    .A2(_1593_),
    .ZN(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5687_ (.I(_0963_),
    .Z(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5688_ (.I(_0958_),
    .Z(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5689_ (.A1(_1595_),
    .A2(_0318_),
    .B1(_3368_),
    .B2(_1596_),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5690_ (.A1(_0963_),
    .A2(_0313_),
    .A3(_0314_),
    .A4(_0959_),
    .ZN(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5691_ (.I(_1599_),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5692_ (.A1(_1597_),
    .A2(_1600_),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5693_ (.A1(_1592_),
    .A2(_1593_),
    .Z(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5694_ (.A1(_1601_),
    .A2(_1602_),
    .ZN(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5695_ (.A1(_1594_),
    .A2(_1603_),
    .ZN(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5696_ (.A1(_0327_),
    .A2(_0972_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5697_ (.A1(_1326_),
    .A2(_1605_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5698_ (.I(_1606_),
    .Z(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5699_ (.A1(_0325_),
    .A2(_0969_),
    .A3(_1607_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5700_ (.A1(_1357_),
    .A2(_1366_),
    .Z(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5701_ (.A1(_1608_),
    .A2(_1610_),
    .ZN(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5702_ (.I(_0326_),
    .Z(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5703_ (.A1(_1612_),
    .A2(_1156_),
    .A3(_1607_),
    .A4(_1610_),
    .Z(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5704_ (.A1(_1604_),
    .A2(_1611_),
    .B(_1613_),
    .ZN(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5705_ (.A1(_1353_),
    .A2(_1354_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5706_ (.A1(_1352_),
    .A2(_1355_),
    .ZN(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5707_ (.A1(_1615_),
    .A2(_1616_),
    .ZN(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5708_ (.A1(_1614_),
    .A2(_1617_),
    .Z(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5709_ (.A1(_0668_),
    .A2(_0342_),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5710_ (.I(_1619_),
    .ZN(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5711_ (.A1(_1614_),
    .A2(_1617_),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5712_ (.A1(_1618_),
    .A2(_1621_),
    .B(_1622_),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5713_ (.A1(_1388_),
    .A2(_1391_),
    .ZN(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5714_ (.A1(_1604_),
    .A2(_1611_),
    .Z(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5715_ (.A1(_0325_),
    .A2(_0969_),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5716_ (.A1(_1607_),
    .A2(_1626_),
    .Z(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5717_ (.A1(_0411_),
    .A2(_0998_),
    .B1(_1000_),
    .B2(_0328_),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5718_ (.A1(_0693_),
    .A2(_3390_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5719_ (.A1(_0917_),
    .A2(_0114_),
    .ZN(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5720_ (.A1(_0065_),
    .A2(_0690_),
    .ZN(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5721_ (.A1(_0694_),
    .A2(_0220_),
    .B1(_0149_),
    .B2(_0687_),
    .ZN(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5722_ (.A1(_1629_),
    .A2(_1630_),
    .B1(_1632_),
    .B2(_1633_),
    .ZN(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5723_ (.A1(_1295_),
    .A2(_1629_),
    .A3(_1339_),
    .ZN(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5724_ (.A1(_1634_),
    .A2(_1635_),
    .ZN(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5725_ (.A1(_1634_),
    .A2(_1635_),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5726_ (.A1(_1607_),
    .A2(_1628_),
    .A3(_1636_),
    .B(_1637_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5727_ (.A1(_1336_),
    .A2(_1343_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5728_ (.A1(_1638_),
    .A2(_1639_),
    .ZN(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5729_ (.A1(_1638_),
    .A2(_1639_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5730_ (.A1(_1627_),
    .A2(_1640_),
    .B(_1641_),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5731_ (.A1(_1335_),
    .A2(_1348_),
    .Z(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5732_ (.A1(_1643_),
    .A2(_1644_),
    .Z(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5733_ (.A1(_1643_),
    .A2(_1644_),
    .Z(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5734_ (.A1(_1625_),
    .A2(_1645_),
    .B(_1646_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5735_ (.A1(_1350_),
    .A2(_1390_),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5736_ (.A1(_1387_),
    .A2(_1648_),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5737_ (.A1(_1618_),
    .A2(_1621_),
    .Z(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5738_ (.I(_1650_),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5739_ (.A1(_1387_),
    .A2(_1648_),
    .Z(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5740_ (.A1(_1647_),
    .A2(_1652_),
    .Z(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5741_ (.A1(_1624_),
    .A2(_1647_),
    .A3(_1649_),
    .B1(_1651_),
    .B2(_1654_),
    .ZN(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5742_ (.A1(_1459_),
    .A2(_1460_),
    .Z(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5743_ (.A1(_1655_),
    .A2(_1656_),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5744_ (.A1(_1655_),
    .A2(_1656_),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5745_ (.A1(_1623_),
    .A2(_1657_),
    .B(_1658_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5746_ (.A1(_1522_),
    .A2(_1524_),
    .Z(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5747_ (.A1(_1659_),
    .A2(_1660_),
    .Z(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5748_ (.A1(_1623_),
    .A2(_1657_),
    .Z(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5749_ (.A1(_1651_),
    .A2(_1654_),
    .ZN(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5750_ (.A1(_1601_),
    .A2(_1602_),
    .Z(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5751_ (.A1(_0392_),
    .A2(_0946_),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5752_ (.A1(_3367_),
    .A2(_1043_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5753_ (.A1(_0948_),
    .A2(_0395_),
    .B1(_0953_),
    .B2(_3367_),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5754_ (.A1(_3297_),
    .A2(_0830_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5755_ (.A1(_1666_),
    .A2(_1667_),
    .B1(_1668_),
    .B2(_1669_),
    .ZN(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5756_ (.A1(_1359_),
    .A2(_1666_),
    .A3(_1591_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5757_ (.A1(_1670_),
    .A2(_1671_),
    .ZN(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5758_ (.A1(_1670_),
    .A2(_1671_),
    .Z(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5759_ (.A1(_0387_),
    .A2(_1596_),
    .A3(_1673_),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5760_ (.A1(_1672_),
    .A2(_1674_),
    .ZN(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5761_ (.A1(_1665_),
    .A2(_1676_),
    .ZN(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5762_ (.A1(_1599_),
    .A2(_1677_),
    .Z(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5763_ (.A1(_1665_),
    .A2(_1676_),
    .Z(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5764_ (.I(_1679_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5765_ (.A1(_1062_),
    .A2(_0420_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5766_ (.A1(_0694_),
    .A2(_0114_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5767_ (.A1(_1068_),
    .A2(_0411_),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5768_ (.A1(_3328_),
    .A2(_1007_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5769_ (.A1(_0281_),
    .A2(_1064_),
    .B1(_0546_),
    .B2(_1068_),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5770_ (.A1(_1682_),
    .A2(_1683_),
    .B1(_1684_),
    .B2(_1685_),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5771_ (.A1(_1338_),
    .A2(_1682_),
    .A3(_1632_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5772_ (.A1(_1687_),
    .A2(_1688_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5773_ (.A1(_1687_),
    .A2(_1688_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5774_ (.A1(_1605_),
    .A2(_1689_),
    .B(_1690_),
    .ZN(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5775_ (.A1(_1606_),
    .A2(_1628_),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5776_ (.A1(_1634_),
    .A2(_1635_),
    .Z(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5777_ (.A1(_1692_),
    .A2(_1693_),
    .Z(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5778_ (.A1(_1691_),
    .A2(_1694_),
    .ZN(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5779_ (.A1(_1691_),
    .A2(_1694_),
    .ZN(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5780_ (.A1(_1681_),
    .A2(_1695_),
    .B(_1696_),
    .ZN(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5781_ (.A1(_1627_),
    .A2(_1640_),
    .Z(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5782_ (.A1(_1698_),
    .A2(_1699_),
    .ZN(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5783_ (.A1(_1698_),
    .A2(_1699_),
    .ZN(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5784_ (.A1(_1680_),
    .A2(_1700_),
    .B(_1701_),
    .ZN(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5785_ (.A1(_1625_),
    .A2(_1645_),
    .Z(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5786_ (.A1(_1702_),
    .A2(_1703_),
    .Z(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5787_ (.A1(_1702_),
    .A2(_1703_),
    .Z(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5788_ (.A1(_1678_),
    .A2(_1704_),
    .B(_1705_),
    .ZN(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5789_ (.A1(_1647_),
    .A2(_1652_),
    .ZN(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5790_ (.A1(_1650_),
    .A2(_1707_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5791_ (.A1(_1650_),
    .A2(_1707_),
    .Z(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5792_ (.A1(_1706_),
    .A2(_1710_),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5793_ (.A1(_1600_),
    .A2(_1602_),
    .A3(_1676_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5794_ (.A1(_1663_),
    .A2(_1706_),
    .A3(_1709_),
    .B1(_1711_),
    .B2(_1712_),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5795_ (.A1(_1662_),
    .A2(_1713_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5796_ (.A1(_1702_),
    .A2(_1703_),
    .A3(_1678_),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5797_ (.A1(_0314_),
    .A2(_0953_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5798_ (.A1(_1589_),
    .A2(_1716_),
    .A3(_1669_),
    .Z(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5799_ (.A1(_0318_),
    .A2(_1043_),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5800_ (.A1(_1716_),
    .A2(_1718_),
    .Z(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5801_ (.A1(_1717_),
    .A2(_1720_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5802_ (.I(_1721_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5803_ (.A1(_0387_),
    .A2(_1596_),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5804_ (.A1(_1723_),
    .A2(_1673_),
    .Z(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5805_ (.A1(_1722_),
    .A2(_1724_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5806_ (.A1(_1721_),
    .A2(_1724_),
    .Z(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5807_ (.A1(_0980_),
    .A2(_0257_),
    .ZN(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5808_ (.A1(_0282_),
    .A2(_1064_),
    .ZN(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5809_ (.A1(_1630_),
    .A2(_1728_),
    .A3(_1684_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5810_ (.I(_1068_),
    .Z(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5811_ (.A1(_1731_),
    .A2(_0351_),
    .A3(_0350_),
    .A4(_1140_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5812_ (.A1(_1729_),
    .A2(_1732_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5813_ (.A1(_1605_),
    .A2(_1687_),
    .A3(_1688_),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5814_ (.A1(_1733_),
    .A2(_1734_),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5815_ (.A1(_1733_),
    .A2(_1734_),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5816_ (.A1(_1727_),
    .A2(_1735_),
    .B(_1736_),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5817_ (.A1(_1691_),
    .A2(_1694_),
    .A3(_1681_),
    .ZN(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5818_ (.A1(_1737_),
    .A2(_1738_),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5819_ (.A1(_1737_),
    .A2(_1738_),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5820_ (.A1(_1726_),
    .A2(_1739_),
    .B(_1740_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5821_ (.A1(_1698_),
    .A2(_1699_),
    .A3(_1679_),
    .Z(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5822_ (.A1(_1742_),
    .A2(_1743_),
    .Z(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5823_ (.A1(_1742_),
    .A2(_1743_),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5824_ (.A1(_1725_),
    .A2(_1744_),
    .B(_1745_),
    .ZN(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5825_ (.A1(_1715_),
    .A2(_1746_),
    .ZN(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5826_ (.A1(_1737_),
    .A2(_1738_),
    .Z(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5827_ (.A1(_1726_),
    .A2(_1748_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5828_ (.A1(_1717_),
    .A2(_1720_),
    .ZN(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5829_ (.A1(_1722_),
    .A2(_1750_),
    .ZN(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5830_ (.A1(_1729_),
    .A2(_1732_),
    .Z(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5831_ (.A1(_1156_),
    .A2(_0190_),
    .A3(_1753_),
    .Z(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5832_ (.A1(_1733_),
    .A2(_1734_),
    .A3(_1727_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5833_ (.A1(_1754_),
    .A2(_1755_),
    .ZN(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5834_ (.A1(_1754_),
    .A2(_1755_),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5835_ (.A1(_1751_),
    .A2(_1756_),
    .B(_1757_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5836_ (.I(_1758_),
    .ZN(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5837_ (.A1(_1749_),
    .A2(_1759_),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5838_ (.A1(_1725_),
    .A2(_1742_),
    .A3(_1743_),
    .Z(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5839_ (.A1(_1760_),
    .A2(_1761_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5840_ (.A1(_1715_),
    .A2(_1746_),
    .Z(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5841_ (.A1(_1726_),
    .A2(_1748_),
    .A3(_1758_),
    .Z(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5842_ (.A1(_1754_),
    .A2(_1755_),
    .A3(_1751_),
    .Z(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5843_ (.A1(_1156_),
    .A2(_0190_),
    .B(_1753_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5844_ (.A1(_1754_),
    .A2(_1767_),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5845_ (.A1(_0476_),
    .A2(_1140_),
    .ZN(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5846_ (.A1(_1683_),
    .A2(_1769_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5847_ (.A1(_1732_),
    .A2(_1770_),
    .ZN(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5848_ (.I(_0980_),
    .Z(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5849_ (.A1(_1772_),
    .A2(_3369_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5850_ (.A1(_1771_),
    .A2(_1773_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5851_ (.A1(_0341_),
    .A2(_1039_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5852_ (.I(_1720_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5853_ (.A1(_1667_),
    .A2(_1776_),
    .B(_1777_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5854_ (.A1(_1768_),
    .A2(_1775_),
    .Z(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5855_ (.A1(_1768_),
    .A2(_1775_),
    .B1(_1778_),
    .B2(_1779_),
    .ZN(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5856_ (.A1(_1765_),
    .A2(_1766_),
    .A3(_1780_),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5857_ (.A1(_1765_),
    .A2(_1766_),
    .A3(_1780_),
    .B1(_1759_),
    .B2(_1749_),
    .ZN(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5858_ (.A1(_1761_),
    .A2(_1782_),
    .Z(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5859_ (.A1(_1766_),
    .A2(_1780_),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5860_ (.A1(_1778_),
    .A2(_1779_),
    .Z(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5861_ (.A1(_1771_),
    .A2(_1773_),
    .Z(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5862_ (.A1(_1731_),
    .A2(_0476_),
    .A3(_1772_),
    .A4(_0342_),
    .Z(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5863_ (.A1(_1787_),
    .A2(_1788_),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5864_ (.A1(_1787_),
    .A2(_1788_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5865_ (.A1(_1718_),
    .A2(_1789_),
    .B(_1790_),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5866_ (.A1(_1786_),
    .A2(_1791_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5867_ (.A1(_1765_),
    .A2(_1784_),
    .A3(_1792_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5868_ (.A1(_1761_),
    .A2(_1781_),
    .B1(_1783_),
    .B2(_1793_),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5869_ (.A1(_1762_),
    .A2(_1715_),
    .A3(_1746_),
    .Z(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5870_ (.A1(_1762_),
    .A2(_1747_),
    .A3(_1764_),
    .B1(_1794_),
    .B2(_1795_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _5871_ (.A1(_1712_),
    .A2(_1706_),
    .A3(_1710_),
    .Z(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5872_ (.A1(_1797_),
    .A2(_1798_),
    .Z(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5873_ (.A1(_1797_),
    .A2(_1798_),
    .Z(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5874_ (.A1(_1747_),
    .A2(_1799_),
    .B(_1800_),
    .ZN(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5875_ (.A1(_1659_),
    .A2(_1660_),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5876_ (.A1(_1662_),
    .A2(_1713_),
    .ZN(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5877_ (.A1(_1714_),
    .A2(_1801_),
    .B(_1802_),
    .C(_1803_),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5878_ (.A1(_1586_),
    .A2(_1661_),
    .A3(_1804_),
    .Z(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5879_ (.A1(_1584_),
    .A2(_1805_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5880_ (.A1(_1470_),
    .A2(_1518_),
    .Z(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5881_ (.A1(_1529_),
    .A2(_1808_),
    .B(_1581_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5882_ (.A1(_1528_),
    .A2(_1582_),
    .ZN(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5883_ (.I(_1526_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5884_ (.A1(_1811_),
    .A2(_0530_),
    .A3(_1578_),
    .ZN(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5885_ (.A1(_1573_),
    .A2(_1577_),
    .B(_1812_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5886_ (.A1(_1534_),
    .A2(_1571_),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5887_ (.A1(_1534_),
    .A2(_1571_),
    .ZN(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5888_ (.A1(_1814_),
    .A2(_1580_),
    .B(_1815_),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5889_ (.I(_0420_),
    .Z(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5890_ (.A1(_1199_),
    .A2(_1817_),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5891_ (.A1(_1561_),
    .A2(_1567_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5892_ (.A1(_1563_),
    .A2(_1820_),
    .ZN(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5893_ (.A1(_1559_),
    .A2(_1569_),
    .Z(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5894_ (.A1(_1559_),
    .A2(_1569_),
    .Z(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5895_ (.A1(_1556_),
    .A2(_1822_),
    .B(_1823_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5896_ (.A1(_1821_),
    .A2(_1824_),
    .Z(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5897_ (.A1(_1819_),
    .A2(_1825_),
    .Z(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5898_ (.A1(_1536_),
    .A2(_1552_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5899_ (.A1(_1553_),
    .A2(_1570_),
    .B(_1827_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5900_ (.A1(_1508_),
    .A2(_1511_),
    .B1(_1560_),
    .B2(_1568_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5901_ (.A1(_1546_),
    .A2(_1549_),
    .ZN(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5902_ (.A1(_1546_),
    .A2(_1549_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5903_ (.A1(_1548_),
    .A2(_1831_),
    .A3(_1832_),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5904_ (.A1(_1545_),
    .A2(_1550_),
    .B(_1833_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5905_ (.A1(_1229_),
    .A2(_0326_),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5906_ (.A1(_0287_),
    .A2(_0959_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5907_ (.A1(_1562_),
    .A2(_1836_),
    .ZN(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5908_ (.A1(_1835_),
    .A2(_1837_),
    .Z(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _5909_ (.A1(_1830_),
    .A2(_1834_),
    .A3(_1838_),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5910_ (.A1(_1537_),
    .A2(_1542_),
    .Z(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5911_ (.A1(_1544_),
    .A2(_1551_),
    .B(_1841_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5912_ (.A1(_1482_),
    .A2(_1000_),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5913_ (.A1(_1241_),
    .A2(_0562_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5914_ (.A1(_0888_),
    .A2(_1482_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5915_ (.A1(_1539_),
    .A2(_1845_),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5916_ (.A1(_1843_),
    .A2(_1844_),
    .B(_1846_),
    .ZN(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5917_ (.A1(_1247_),
    .A2(_1486_),
    .B1(_1437_),
    .B2(_1222_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5918_ (.A1(_1221_),
    .A2(_0075_),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5919_ (.A1(_1549_),
    .A2(_1849_),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5920_ (.A1(_1848_),
    .A2(_1850_),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5921_ (.A1(_1480_),
    .A2(_1843_),
    .B1(_1541_),
    .B2(_1538_),
    .ZN(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5922_ (.A1(_1852_),
    .A2(_1853_),
    .Z(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5923_ (.A1(_1832_),
    .A2(_1854_),
    .ZN(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5924_ (.A1(_1847_),
    .A2(_1855_),
    .Z(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5925_ (.A1(_1842_),
    .A2(_1856_),
    .Z(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5926_ (.A1(_1839_),
    .A2(_1857_),
    .Z(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5927_ (.A1(_1828_),
    .A2(_1858_),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5928_ (.A1(_1826_),
    .A2(_1859_),
    .Z(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5929_ (.A1(_1816_),
    .A2(_1860_),
    .Z(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5930_ (.A1(_1813_),
    .A2(_1861_),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5931_ (.A1(_1809_),
    .A2(_1810_),
    .B(_1863_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5932_ (.A1(_1809_),
    .A2(_1810_),
    .A3(_1863_),
    .Z(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5933_ (.A1(_1864_),
    .A2(_1865_),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5934_ (.A1(_1806_),
    .A2(_1866_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5935_ (.A1(_1274_),
    .A2(_1867_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5936_ (.A1(_3294_),
    .A2(_1266_),
    .B(_1270_),
    .C(_1868_),
    .ZN(net19));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5937_ (.A1(_0383_),
    .A2(_0514_),
    .A3(_0519_),
    .Z(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5938_ (.A1(_0303_),
    .A2(_0582_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5939_ (.A1(_0303_),
    .A2(_0524_),
    .A3(_0582_),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5940_ (.A1(_0529_),
    .A2(_0580_),
    .ZN(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5941_ (.A1(_0244_),
    .A2(_0301_),
    .B1(_0529_),
    .B2(_0580_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5942_ (.A1(_1873_),
    .A2(_1874_),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5943_ (.A1(_1869_),
    .A2(_1870_),
    .B(_1871_),
    .C(_1875_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5944_ (.I(_2909_),
    .Z(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5945_ (.A1(_1877_),
    .A2(_1817_),
    .A3(_0541_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5946_ (.A1(_0537_),
    .A2(_0540_),
    .B(_1878_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5947_ (.A1(_0544_),
    .A2(_0576_),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5948_ (.A1(_0542_),
    .A2(_0577_),
    .B(_1880_),
    .ZN(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5949_ (.A1(_0559_),
    .A2(_0574_),
    .ZN(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5950_ (.A1(_0557_),
    .A2(_0575_),
    .B(_1882_),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5951_ (.A1(_0566_),
    .A2(_0573_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5952_ (.A1(_0075_),
    .A2(_2809_),
    .ZN(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5953_ (.A1(_0561_),
    .A2(_1301_),
    .Z(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5954_ (.A1(_1886_),
    .A2(_1887_),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5955_ (.A1(_0565_),
    .A2(_1888_),
    .Z(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5956_ (.A1(_0568_),
    .A2(_1889_),
    .ZN(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5957_ (.A1(_0564_),
    .A2(_1890_),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5958_ (.A1(_1885_),
    .A2(_1891_),
    .Z(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5959_ (.A1(_0569_),
    .A2(_0571_),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5960_ (.A1(_0273_),
    .A2(_0572_),
    .ZN(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5961_ (.A1(_1893_),
    .A2(_1895_),
    .ZN(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5962_ (.I(_0287_),
    .Z(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5963_ (.I(_3251_),
    .Z(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5964_ (.A1(_1897_),
    .A2(_0317_),
    .B1(_1898_),
    .B2(_1564_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5965_ (.A1(_1897_),
    .A2(_3251_),
    .ZN(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5966_ (.A1(_0290_),
    .A2(_1900_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5967_ (.A1(_1899_),
    .A2(_1901_),
    .ZN(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5968_ (.A1(_1896_),
    .A2(_1902_),
    .Z(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5969_ (.A1(_1892_),
    .A2(_1903_),
    .Z(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5970_ (.A1(_1884_),
    .A2(_1904_),
    .Z(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5971_ (.A1(_0551_),
    .A2(_0555_),
    .Z(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5972_ (.A1(_0545_),
    .A2(_0556_),
    .B(_1907_),
    .ZN(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5973_ (.A1(_0290_),
    .A2(_0553_),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5974_ (.A1(_0552_),
    .A2(_0554_),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5975_ (.A1(_1909_),
    .A2(_1910_),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5976_ (.A1(_1908_),
    .A2(_1911_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5977_ (.A1(_1612_),
    .A2(_2908_),
    .ZN(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5978_ (.A1(_1912_),
    .A2(_1913_),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5979_ (.A1(_1906_),
    .A2(_1914_),
    .Z(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5980_ (.A1(_1881_),
    .A2(_1915_),
    .Z(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5981_ (.A1(_1879_),
    .A2(_1917_),
    .ZN(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5982_ (.A1(_0534_),
    .A2(_0578_),
    .Z(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5983_ (.A1(_0532_),
    .A2(_0579_),
    .B(_1919_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5984_ (.A1(_1918_),
    .A2(_1920_),
    .Z(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5985_ (.A1(_1876_),
    .A2(_1921_),
    .Z(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5986_ (.I(net16),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5987_ (.A1(_1923_),
    .A2(_1271_),
    .ZN(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5988_ (.I(_1924_),
    .Z(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5989_ (.A1(_1876_),
    .A2(_1921_),
    .B(_1925_),
    .ZN(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5990_ (.A1(_1922_),
    .A2(_1926_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5991_ (.A1(_0696_),
    .A2(_1928_),
    .ZN(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5992_ (.A1(_3220_),
    .A2(_3287_),
    .Z(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5993_ (.A1(_3220_),
    .A2(_3218_),
    .A3(_3287_),
    .Z(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5994_ (.A1(_3224_),
    .A2(_3286_),
    .Z(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5995_ (.A1(_3224_),
    .A2(_3286_),
    .Z(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5996_ (.A1(_2981_),
    .A2(_1932_),
    .B(_1933_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5997_ (.A1(_3215_),
    .A2(_1930_),
    .B(_1931_),
    .C(_1934_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5998_ (.A1(_1877_),
    .A2(_1208_),
    .A3(_3238_),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5999_ (.A1(_3234_),
    .A2(_3237_),
    .B(_1936_),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6000_ (.A1(_3241_),
    .A2(_3283_),
    .ZN(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6001_ (.A1(_3239_),
    .A2(_3284_),
    .B(_1939_),
    .ZN(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6002_ (.A1(_3259_),
    .A2(_3281_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6003_ (.A1(_3257_),
    .A2(_3282_),
    .B(_1941_),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6004_ (.A1(_3268_),
    .A2(_3280_),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6005_ (.A1(_3269_),
    .A2(_3244_),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6006_ (.A1(_3263_),
    .A2(_3274_),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6007_ (.A1(_1944_),
    .A2(_1945_),
    .Z(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6008_ (.A1(_3267_),
    .A2(_1946_),
    .Z(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6009_ (.A1(_3275_),
    .A2(_1947_),
    .ZN(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6010_ (.A1(_3266_),
    .A2(_1948_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6011_ (.A1(_1943_),
    .A2(_1950_),
    .Z(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6012_ (.A1(_3276_),
    .A2(_3278_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6013_ (.A1(_2970_),
    .A2(_3279_),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6014_ (.A1(_1952_),
    .A2(_1953_),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6015_ (.I(_2938_),
    .Z(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6016_ (.A1(_1955_),
    .A2(_0317_),
    .B1(_1378_),
    .B2(_1898_),
    .ZN(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6017_ (.A1(_1955_),
    .A2(_1898_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6018_ (.A1(_2946_),
    .A2(_1957_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6019_ (.A1(_1956_),
    .A2(_1958_),
    .ZN(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6020_ (.A1(_1954_),
    .A2(_1959_),
    .Z(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6021_ (.A1(_1951_),
    .A2(_1961_),
    .Z(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6022_ (.A1(_1942_),
    .A2(_1962_),
    .Z(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6023_ (.A1(_3250_),
    .A2(_3255_),
    .Z(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6024_ (.A1(_3242_),
    .A2(_3256_),
    .B(_1964_),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6025_ (.A1(_2946_),
    .A2(_3253_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6026_ (.A1(_3252_),
    .A2(_3254_),
    .ZN(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6027_ (.A1(_1966_),
    .A2(_1967_),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6028_ (.A1(_1965_),
    .A2(_1968_),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6029_ (.A1(_0979_),
    .A2(_2908_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6030_ (.A1(_1969_),
    .A2(_1970_),
    .Z(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6031_ (.A1(_1963_),
    .A2(_1972_),
    .Z(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6032_ (.A1(_1940_),
    .A2(_1973_),
    .Z(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6033_ (.A1(_1937_),
    .A2(_1974_),
    .Z(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6034_ (.A1(_3231_),
    .A2(_3285_),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6035_ (.A1(_3231_),
    .A2(_3285_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6036_ (.A1(_3228_),
    .A2(_1976_),
    .B(_1977_),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6037_ (.A1(_1975_),
    .A2(_1978_),
    .ZN(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6038_ (.A1(_1935_),
    .A2(_1979_),
    .Z(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6039_ (.A1(_1923_),
    .A2(_0674_),
    .ZN(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6040_ (.A1(_1935_),
    .A2(_1979_),
    .B(_1981_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6041_ (.A1(_1526_),
    .A2(_1208_),
    .A3(_1216_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6042_ (.A1(_1211_),
    .A2(_1215_),
    .B(_1984_),
    .ZN(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6043_ (.A1(_1219_),
    .A2(_1260_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6044_ (.A1(_1217_),
    .A2(_1261_),
    .B(_1986_),
    .ZN(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6045_ (.A1(_1238_),
    .A2(_1258_),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6046_ (.A1(_1236_),
    .A2(_1259_),
    .B(_1988_),
    .ZN(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6047_ (.A1(_1245_),
    .A2(_1256_),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6048_ (.A1(_1221_),
    .A2(_3269_),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6049_ (.A1(_1250_),
    .A2(_3263_),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6050_ (.A1(_1991_),
    .A2(_1992_),
    .Z(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6051_ (.A1(_1244_),
    .A2(_1994_),
    .Z(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6052_ (.A1(_1251_),
    .A2(_1995_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6053_ (.A1(_1243_),
    .A2(_1996_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6054_ (.A1(_1990_),
    .A2(_1997_),
    .Z(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6055_ (.A1(_1252_),
    .A2(_1254_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6056_ (.A1(_0857_),
    .A2(_1255_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6057_ (.A1(_1999_),
    .A2(_2000_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6058_ (.I(_1955_),
    .Z(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6059_ (.I(_1378_),
    .Z(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6060_ (.I(_1229_),
    .Z(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6061_ (.A1(_1595_),
    .A2(_2002_),
    .B1(_2003_),
    .B2(_2005_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6062_ (.A1(_2005_),
    .A2(_1955_),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6063_ (.A1(_0834_),
    .A2(_2007_),
    .ZN(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6064_ (.A1(_2006_),
    .A2(_2008_),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6065_ (.A1(_2001_),
    .A2(_2009_),
    .Z(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6066_ (.A1(_1998_),
    .A2(_2010_),
    .Z(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6067_ (.A1(_1989_),
    .A2(_2011_),
    .Z(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6068_ (.A1(_1227_),
    .A2(_1233_),
    .Z(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6069_ (.A1(_1220_),
    .A2(_1234_),
    .B(_2013_),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6070_ (.A1(_0834_),
    .A2(_1231_),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6071_ (.A1(_1230_),
    .A2(_1232_),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6072_ (.A1(_2016_),
    .A2(_2017_),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6073_ (.A1(_2014_),
    .A2(_2018_),
    .Z(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6074_ (.A1(_2014_),
    .A2(_2018_),
    .ZN(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6075_ (.A1(_2019_),
    .A2(_2020_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6076_ (.A1(_0669_),
    .A2(_0979_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6077_ (.A1(_2021_),
    .A2(_2022_),
    .Z(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6078_ (.A1(_2012_),
    .A2(_2023_),
    .Z(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6079_ (.A1(_1987_),
    .A2(_2024_),
    .Z(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6080_ (.A1(_1985_),
    .A2(_2025_),
    .Z(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6081_ (.A1(_1207_),
    .A2(_1262_),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6082_ (.A1(_1207_),
    .A2(_1262_),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6083_ (.A1(_1204_),
    .A2(_2028_),
    .B(_2029_),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6084_ (.A1(_2027_),
    .A2(_2030_),
    .Z(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6085_ (.A1(_1198_),
    .A2(_1263_),
    .Z(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6086_ (.A1(_0945_),
    .A2(_2032_),
    .Z(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6087_ (.A1(_1198_),
    .A2(_1263_),
    .Z(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6088_ (.A1(_1195_),
    .A2(_2033_),
    .B(_2034_),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6089_ (.A1(_2031_),
    .A2(_2035_),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6090_ (.A1(_2027_),
    .A2(_2030_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6091_ (.A1(_1194_),
    .A2(_1264_),
    .Z(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6092_ (.A1(_1194_),
    .A2(_1193_),
    .A3(_1264_),
    .Z(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6093_ (.A1(_0945_),
    .A2(_2034_),
    .B(_2032_),
    .ZN(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6094_ (.A1(_1188_),
    .A2(_2039_),
    .B(_2040_),
    .C(_2041_),
    .ZN(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6095_ (.A1(_1923_),
    .A2(_1271_),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6096_ (.I(_2043_),
    .Z(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6097_ (.A1(_2038_),
    .A2(_2042_),
    .B(_2044_),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6098_ (.A1(_1980_),
    .A2(_1983_),
    .B1(_2036_),
    .B2(_2045_),
    .ZN(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6099_ (.A1(_1811_),
    .A2(_1817_),
    .A3(_1825_),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6100_ (.A1(_1821_),
    .A2(_1824_),
    .B(_2047_),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6101_ (.A1(_1828_),
    .A2(_1858_),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6102_ (.A1(_1826_),
    .A2(_1859_),
    .B(_2050_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6103_ (.I(_1842_),
    .ZN(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6104_ (.A1(_2052_),
    .A2(_1856_),
    .ZN(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6105_ (.A1(_1839_),
    .A2(_1857_),
    .B(_2053_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6106_ (.I(_1854_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6107_ (.A1(_1852_),
    .A2(_1853_),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6108_ (.A1(_1832_),
    .A2(_2055_),
    .B(_2056_),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6109_ (.I(_1897_),
    .Z(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6110_ (.A1(_1595_),
    .A2(_2058_),
    .B1(_2005_),
    .B2(_1564_),
    .ZN(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6111_ (.A1(_1897_),
    .A2(_1229_),
    .ZN(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6112_ (.A1(_1562_),
    .A2(_2061_),
    .ZN(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6113_ (.A1(_2060_),
    .A2(_2062_),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6114_ (.A1(_2057_),
    .A2(_2063_),
    .Z(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6115_ (.A1(_1847_),
    .A2(_1855_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6116_ (.A1(_1250_),
    .A2(_0562_),
    .ZN(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6117_ (.A1(_1849_),
    .A2(_2066_),
    .Z(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6118_ (.A1(_1846_),
    .A2(_2067_),
    .Z(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6119_ (.A1(_1850_),
    .A2(_2068_),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6120_ (.A1(_1845_),
    .A2(_2069_),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6121_ (.A1(_2065_),
    .A2(_2071_),
    .Z(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6122_ (.A1(_2064_),
    .A2(_2072_),
    .Z(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6123_ (.A1(_2054_),
    .A2(_2073_),
    .Z(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6124_ (.A1(_1834_),
    .A2(_1838_),
    .Z(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6125_ (.A1(_1834_),
    .A2(_1838_),
    .Z(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6126_ (.A1(_1830_),
    .A2(_2075_),
    .B(_2076_),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6127_ (.A1(_1562_),
    .A2(_1836_),
    .ZN(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6128_ (.A1(_1835_),
    .A2(_1837_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6129_ (.A1(_2078_),
    .A2(_2079_),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6130_ (.A1(_2077_),
    .A2(_2080_),
    .Z(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6131_ (.A1(_2077_),
    .A2(_2080_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6132_ (.A1(_2082_),
    .A2(_2083_),
    .ZN(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6133_ (.A1(_0669_),
    .A2(_1612_),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6134_ (.A1(_2084_),
    .A2(_2085_),
    .Z(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6135_ (.A1(_2074_),
    .A2(_2086_),
    .Z(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6136_ (.A1(_2051_),
    .A2(_2087_),
    .Z(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6137_ (.A1(_2049_),
    .A2(_2088_),
    .ZN(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6138_ (.A1(_1816_),
    .A2(_1860_),
    .ZN(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6139_ (.A1(_1813_),
    .A2(_1861_),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6140_ (.A1(_2090_),
    .A2(_2091_),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6141_ (.A1(_2089_),
    .A2(_2093_),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6142_ (.A1(_1586_),
    .A2(_1661_),
    .A3(_1804_),
    .A4(_1866_),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6143_ (.I(_1865_),
    .ZN(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6144_ (.A1(_1584_),
    .A2(_1864_),
    .B(_2096_),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6145_ (.A1(_2095_),
    .A2(_2097_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6146_ (.A1(_2094_),
    .A2(_2098_),
    .Z(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6147_ (.A1(_1274_),
    .A2(_2099_),
    .ZN(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6148_ (.A1(_1929_),
    .A2(_2046_),
    .B(_1270_),
    .C(_2100_),
    .ZN(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6149_ (.I(_0685_),
    .Z(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6150_ (.I(_2101_),
    .Z(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6151_ (.A1(_2051_),
    .A2(_2087_),
    .ZN(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6152_ (.A1(_2049_),
    .A2(_2088_),
    .ZN(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6153_ (.A1(_2084_),
    .A2(_2085_),
    .B(_2082_),
    .ZN(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6154_ (.A1(_2054_),
    .A2(_2073_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6155_ (.A1(_2074_),
    .A2(_2086_),
    .ZN(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6156_ (.A1(_2107_),
    .A2(_2108_),
    .ZN(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6157_ (.A1(_2064_),
    .A2(_2072_),
    .ZN(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6158_ (.A1(_2065_),
    .A2(_2071_),
    .B(_2110_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6159_ (.A1(_1845_),
    .A2(_2069_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6160_ (.I(_1482_),
    .Z(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6161_ (.I(_0824_),
    .Z(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6162_ (.A1(_2114_),
    .A2(_2115_),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6163_ (.I(_2115_),
    .Z(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6164_ (.I(_1486_),
    .Z(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6165_ (.I(_0562_),
    .Z(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6166_ (.I(_1223_),
    .Z(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6167_ (.A1(_2119_),
    .A2(_2120_),
    .ZN(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6168_ (.A1(_2117_),
    .A2(_2118_),
    .B(_2121_),
    .ZN(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6169_ (.A1(_2116_),
    .A2(_2122_),
    .Z(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6170_ (.A1(_2112_),
    .A2(_2123_),
    .Z(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6171_ (.A1(_1846_),
    .A2(_2067_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6172_ (.A1(_1850_),
    .A2(_2068_),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6173_ (.A1(_2126_),
    .A2(_2127_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6174_ (.A1(_2061_),
    .A2(_2128_),
    .Z(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6175_ (.A1(_2125_),
    .A2(_2129_),
    .Z(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6176_ (.I(_1564_),
    .Z(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6177_ (.A1(_2131_),
    .A2(_0670_),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6178_ (.A1(_2057_),
    .A2(_2062_),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6179_ (.A1(_2060_),
    .A2(_2133_),
    .ZN(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6180_ (.A1(_2132_),
    .A2(_2134_),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6181_ (.A1(_2111_),
    .A2(_2130_),
    .A3(_2136_),
    .Z(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6182_ (.A1(_2106_),
    .A2(_2109_),
    .A3(_2137_),
    .Z(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6183_ (.A1(_2104_),
    .A2(_2105_),
    .B(_2138_),
    .ZN(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6184_ (.A1(_2104_),
    .A2(_2105_),
    .A3(_2138_),
    .Z(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6185_ (.A1(_2139_),
    .A2(_2140_),
    .ZN(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6186_ (.A1(_2090_),
    .A2(_2091_),
    .B(_2089_),
    .ZN(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6187_ (.A1(_2094_),
    .A2(_2098_),
    .B(_2142_),
    .ZN(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6188_ (.A1(_2141_),
    .A2(_2143_),
    .Z(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6189_ (.I(_3290_),
    .Z(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6190_ (.I(_2145_),
    .Z(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6191_ (.A1(_1940_),
    .A2(_1973_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6192_ (.A1(_1937_),
    .A2(_1974_),
    .ZN(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6193_ (.A1(_1965_),
    .A2(_1968_),
    .Z(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6194_ (.A1(_1969_),
    .A2(_1970_),
    .B(_2150_),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6195_ (.A1(_1942_),
    .A2(_1962_),
    .ZN(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6196_ (.A1(_1963_),
    .A2(_1972_),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6197_ (.A1(_2152_),
    .A2(_2153_),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6198_ (.A1(_1951_),
    .A2(_1961_),
    .ZN(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6199_ (.A1(_1943_),
    .A2(_1950_),
    .B(_2155_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6200_ (.A1(_3266_),
    .A2(_1948_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6201_ (.A1(_1239_),
    .A2(_3243_),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6202_ (.I(_3270_),
    .Z(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6203_ (.A1(_3264_),
    .A2(_3245_),
    .ZN(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6204_ (.A1(_3243_),
    .A2(_2160_),
    .B(_2161_),
    .ZN(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6205_ (.A1(_2159_),
    .A2(_2162_),
    .Z(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6206_ (.A1(_2158_),
    .A2(_2163_),
    .Z(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6207_ (.A1(_3267_),
    .A2(_1946_),
    .ZN(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6208_ (.A1(_3275_),
    .A2(_1947_),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6209_ (.A1(_2165_),
    .A2(_2166_),
    .ZN(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6210_ (.A1(_1957_),
    .A2(_2167_),
    .Z(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6211_ (.A1(_2164_),
    .A2(_2169_),
    .Z(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6212_ (.A1(_2156_),
    .A2(_2170_),
    .Z(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6213_ (.I(_2907_),
    .Z(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6214_ (.A1(_2003_),
    .A2(_2172_),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6215_ (.I(_1956_),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6216_ (.A1(_1954_),
    .A2(_1958_),
    .B(_2174_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6217_ (.A1(_2173_),
    .A2(_2175_),
    .Z(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6218_ (.A1(_2171_),
    .A2(_2176_),
    .ZN(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6219_ (.A1(_2151_),
    .A2(_2154_),
    .A3(_2177_),
    .Z(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6220_ (.A1(_2148_),
    .A2(_2149_),
    .B(_2178_),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6221_ (.A1(_2148_),
    .A2(_2149_),
    .A3(_2178_),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6222_ (.I(_2181_),
    .ZN(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6223_ (.A1(_2180_),
    .A2(_2182_),
    .Z(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6224_ (.A1(_1975_),
    .A2(_1978_),
    .ZN(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6225_ (.A1(_2184_),
    .A2(_1980_),
    .ZN(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6226_ (.A1(_2183_),
    .A2(_2185_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6227_ (.A1(_2147_),
    .A2(_2186_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6228_ (.A1(_1918_),
    .A2(_1920_),
    .ZN(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6229_ (.A1(_1908_),
    .A2(_1911_),
    .Z(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6230_ (.A1(_1912_),
    .A2(_1913_),
    .B(_2189_),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6231_ (.A1(_1884_),
    .A2(_1904_),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6232_ (.A1(_1906_),
    .A2(_1914_),
    .ZN(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6233_ (.A1(_2192_),
    .A2(_2193_),
    .ZN(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6234_ (.A1(_1892_),
    .A2(_1903_),
    .ZN(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6235_ (.A1(_1885_),
    .A2(_1891_),
    .B(_2195_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6236_ (.A1(_0564_),
    .A2(_1890_),
    .ZN(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6237_ (.I(_3243_),
    .Z(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6238_ (.A1(_2114_),
    .A2(_2198_),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6239_ (.I(_3245_),
    .Z(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6240_ (.A1(_2119_),
    .A2(_2200_),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6241_ (.A1(_2118_),
    .A2(_2198_),
    .B(_2202_),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6242_ (.A1(_2199_),
    .A2(_2203_),
    .Z(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6243_ (.A1(_2197_),
    .A2(_2204_),
    .Z(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6244_ (.A1(_0565_),
    .A2(_1888_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6245_ (.A1(_0568_),
    .A2(_1889_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6246_ (.A1(_2206_),
    .A2(_2207_),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6247_ (.A1(_1900_),
    .A2(_2208_),
    .Z(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6248_ (.A1(_2205_),
    .A2(_2209_),
    .Z(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6249_ (.A1(_2196_),
    .A2(_2210_),
    .Z(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6250_ (.A1(_2131_),
    .A2(_2172_),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6251_ (.I(_1899_),
    .ZN(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6252_ (.A1(_1896_),
    .A2(_1901_),
    .B(_2214_),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6253_ (.A1(_2213_),
    .A2(_2215_),
    .Z(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6254_ (.A1(_2211_),
    .A2(_2216_),
    .ZN(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6255_ (.A1(_2191_),
    .A2(_2194_),
    .A3(_2217_),
    .Z(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6256_ (.A1(_1881_),
    .A2(_1915_),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6257_ (.A1(_1879_),
    .A2(_1917_),
    .ZN(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6258_ (.A1(_2219_),
    .A2(_2220_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6259_ (.A1(_2218_),
    .A2(_2221_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6260_ (.A1(_2188_),
    .A2(_1922_),
    .B(_2222_),
    .ZN(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6261_ (.I(_0674_),
    .Z(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6262_ (.A1(_3295_),
    .A2(_2225_),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6263_ (.A1(_2188_),
    .A2(_1922_),
    .A3(_2222_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6264_ (.A1(_2226_),
    .A2(_2227_),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6265_ (.A1(_2027_),
    .A2(_2030_),
    .Z(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6266_ (.A1(_2031_),
    .A2(_2035_),
    .B(_2229_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6267_ (.A1(_2021_),
    .A2(_2022_),
    .B(_2019_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6268_ (.A1(_1989_),
    .A2(_2011_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6269_ (.A1(_2012_),
    .A2(_2023_),
    .ZN(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6270_ (.A1(_2232_),
    .A2(_2233_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6271_ (.A1(_1998_),
    .A2(_2010_),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6272_ (.A1(_1990_),
    .A2(_1997_),
    .B(_2236_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6273_ (.A1(_1243_),
    .A2(_1996_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6274_ (.A1(_2115_),
    .A2(_1239_),
    .ZN(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6275_ (.I(_3264_),
    .Z(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6276_ (.A1(_1223_),
    .A2(_2240_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6277_ (.A1(_2115_),
    .A2(_2160_),
    .B(_2241_),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6278_ (.A1(_2239_),
    .A2(_2242_),
    .Z(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6279_ (.A1(_2238_),
    .A2(_2243_),
    .Z(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6280_ (.A1(_1244_),
    .A2(_1994_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6281_ (.A1(_1251_),
    .A2(_1995_),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6282_ (.A1(_2246_),
    .A2(_2247_),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6283_ (.A1(_2007_),
    .A2(_2248_),
    .Z(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6284_ (.A1(_2244_),
    .A2(_2249_),
    .Z(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6285_ (.A1(_2237_),
    .A2(_2250_),
    .Z(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6286_ (.A1(_1200_),
    .A2(_2003_),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6287_ (.I(_2006_),
    .ZN(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6288_ (.A1(_2001_),
    .A2(_2008_),
    .B(_2253_),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6289_ (.A1(_2252_),
    .A2(_2254_),
    .Z(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6290_ (.A1(_2251_),
    .A2(_2255_),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6291_ (.A1(_2231_),
    .A2(_2235_),
    .A3(_2257_),
    .Z(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6292_ (.A1(_1987_),
    .A2(_2024_),
    .ZN(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6293_ (.A1(_1985_),
    .A2(_2025_),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6294_ (.A1(_2259_),
    .A2(_2260_),
    .ZN(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6295_ (.A1(_2258_),
    .A2(_2261_),
    .Z(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6296_ (.A1(_2230_),
    .A2(_2262_),
    .Z(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6297_ (.I(_0685_),
    .Z(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6298_ (.A1(_2224_),
    .A2(_2228_),
    .B1(_2263_),
    .B2(_0585_),
    .C(_2264_),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6299_ (.I(_1269_),
    .Z(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6300_ (.A1(_2103_),
    .A2(_2144_),
    .B1(_2187_),
    .B2(_2265_),
    .C(_2266_),
    .ZN(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6301_ (.I(_0696_),
    .Z(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6302_ (.A1(_2131_),
    .A2(_1811_),
    .A3(_2134_),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6303_ (.A1(_2111_),
    .A2(_2130_),
    .ZN(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6304_ (.A1(_2111_),
    .A2(_2130_),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6305_ (.A1(_2270_),
    .A2(_2136_),
    .B(_2271_),
    .ZN(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6306_ (.A1(_2126_),
    .A2(_2127_),
    .B(_2061_),
    .ZN(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6307_ (.A1(_2058_),
    .A2(_0670_),
    .Z(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6308_ (.A1(_1526_),
    .A2(_2273_),
    .ZN(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6309_ (.A1(_2273_),
    .A2(_2274_),
    .B(_2275_),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6310_ (.A1(_1845_),
    .A2(_2069_),
    .A3(_2123_),
    .B1(_2125_),
    .B2(_2129_),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6311_ (.I(_2114_),
    .ZN(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6312_ (.A1(_2279_),
    .A2(_2066_),
    .ZN(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6313_ (.A1(_2279_),
    .A2(_2118_),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6314_ (.A1(_2117_),
    .A2(_2119_),
    .A3(_2281_),
    .ZN(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6315_ (.A1(_2120_),
    .A2(_2280_),
    .A3(_2282_),
    .ZN(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6316_ (.A1(_2278_),
    .A2(_2283_),
    .Z(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6317_ (.A1(_2276_),
    .A2(_2284_),
    .Z(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6318_ (.A1(_2272_),
    .A2(_2285_),
    .Z(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6319_ (.A1(_2269_),
    .A2(_2286_),
    .Z(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6320_ (.I(_2109_),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6321_ (.A1(_2289_),
    .A2(_2137_),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6322_ (.A1(_2289_),
    .A2(_2137_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6323_ (.A1(_2106_),
    .A2(_2290_),
    .B(_2291_),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6324_ (.A1(_2287_),
    .A2(_2292_),
    .Z(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6325_ (.A1(_2094_),
    .A2(_2141_),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6326_ (.A1(_2095_),
    .A2(_2097_),
    .B(_2294_),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6327_ (.A1(_2142_),
    .A2(_2139_),
    .ZN(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6328_ (.A1(_2140_),
    .A2(_2296_),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6329_ (.A1(_2293_),
    .A2(_2295_),
    .A3(_2297_),
    .Z(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6330_ (.A1(_2295_),
    .A2(_2297_),
    .B(_2293_),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6331_ (.A1(_2298_),
    .A2(_2300_),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6332_ (.A1(_2213_),
    .A2(_2215_),
    .ZN(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6333_ (.A1(_2196_),
    .A2(_2210_),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6334_ (.A1(_2211_),
    .A2(_2216_),
    .ZN(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6335_ (.A1(_2303_),
    .A2(_2304_),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6336_ (.A1(_2206_),
    .A2(_2207_),
    .B(_1900_),
    .ZN(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6337_ (.A1(_2058_),
    .A2(_2172_),
    .Z(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6338_ (.A1(_2172_),
    .A2(_2306_),
    .ZN(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6339_ (.A1(_2306_),
    .A2(_2307_),
    .B(_2308_),
    .ZN(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6340_ (.A1(_0564_),
    .A2(_1890_),
    .A3(_2204_),
    .B1(_2205_),
    .B2(_2209_),
    .ZN(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6341_ (.A1(_1887_),
    .A2(_2281_),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6342_ (.A1(_2114_),
    .A2(_1887_),
    .B(_2312_),
    .C(_2200_),
    .ZN(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6343_ (.A1(_2311_),
    .A2(_2313_),
    .Z(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6344_ (.A1(_2309_),
    .A2(_2314_),
    .Z(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6345_ (.A1(_2305_),
    .A2(_2315_),
    .Z(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6346_ (.A1(_2302_),
    .A2(_2316_),
    .ZN(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6347_ (.I(_2194_),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6348_ (.A1(_2318_),
    .A2(_2217_),
    .ZN(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6349_ (.A1(_2318_),
    .A2(_2217_),
    .ZN(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6350_ (.A1(_2191_),
    .A2(_2319_),
    .B(_2320_),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6351_ (.A1(_2317_),
    .A2(_2322_),
    .Z(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6352_ (.A1(_0303_),
    .A2(_0582_),
    .Z(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6353_ (.A1(_0302_),
    .A2(_0524_),
    .A3(_0581_),
    .Z(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6354_ (.A1(_1873_),
    .A2(_1874_),
    .Z(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6355_ (.A1(_0520_),
    .A2(_2324_),
    .B(_2325_),
    .C(_2326_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6356_ (.A1(_1921_),
    .A2(_2222_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6357_ (.A1(_2219_),
    .A2(_2220_),
    .B(_2218_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6358_ (.A1(_2219_),
    .A2(_2220_),
    .A3(_2218_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6359_ (.A1(_2188_),
    .A2(_2329_),
    .B(_2330_),
    .ZN(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6360_ (.A1(_2327_),
    .A2(_2328_),
    .B(_2331_),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6361_ (.A1(_2323_),
    .A2(_2333_),
    .ZN(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6362_ (.A1(_2323_),
    .A2(_2333_),
    .Z(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6363_ (.A1(_1925_),
    .A2(_2334_),
    .A3(_2335_),
    .ZN(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6364_ (.A1(_2252_),
    .A2(_2254_),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6365_ (.A1(_2237_),
    .A2(_2250_),
    .ZN(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6366_ (.A1(_2251_),
    .A2(_2255_),
    .ZN(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6367_ (.A1(_2338_),
    .A2(_2339_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6368_ (.A1(_2246_),
    .A2(_2247_),
    .B(_2007_),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6369_ (.A1(_1200_),
    .A2(_2341_),
    .Z(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6370_ (.A1(_0670_),
    .A2(_2002_),
    .B(_2341_),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6371_ (.A1(_2342_),
    .A2(_2344_),
    .Z(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6372_ (.A1(_1243_),
    .A2(_1996_),
    .A3(_2243_),
    .B1(_2244_),
    .B2(_2249_),
    .ZN(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6373_ (.I(_1239_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6374_ (.A1(_2347_),
    .A2(_1992_),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6375_ (.A1(_2347_),
    .A2(_2160_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6376_ (.A1(_2117_),
    .A2(_2240_),
    .A3(_2349_),
    .ZN(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6377_ (.A1(_2120_),
    .A2(_2348_),
    .A3(_2350_),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6378_ (.A1(_2346_),
    .A2(_2351_),
    .Z(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6379_ (.A1(_2345_),
    .A2(_2352_),
    .Z(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6380_ (.A1(_2340_),
    .A2(_2353_),
    .Z(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6381_ (.A1(_2337_),
    .A2(_2355_),
    .ZN(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6382_ (.I(_2235_),
    .ZN(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6383_ (.A1(_2357_),
    .A2(_2257_),
    .ZN(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6384_ (.A1(_2357_),
    .A2(_2257_),
    .ZN(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6385_ (.A1(_2231_),
    .A2(_2358_),
    .B(_2359_),
    .ZN(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6386_ (.A1(_2356_),
    .A2(_2360_),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6387_ (.A1(_2259_),
    .A2(_2260_),
    .B(_2258_),
    .ZN(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6388_ (.A1(_2259_),
    .A2(_2260_),
    .A3(_2258_),
    .ZN(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6389_ (.A1(_2229_),
    .A2(_2362_),
    .B(_2363_),
    .ZN(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6390_ (.A1(_2038_),
    .A2(_2042_),
    .A3(_2262_),
    .B(_2364_),
    .ZN(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6391_ (.A1(_2361_),
    .A2(_2366_),
    .Z(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6392_ (.I(_0584_),
    .Z(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6393_ (.A1(_2361_),
    .A2(_2366_),
    .B(_2368_),
    .ZN(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6394_ (.A1(_2367_),
    .A2(_2369_),
    .Z(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6395_ (.A1(_2173_),
    .A2(_2175_),
    .Z(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6396_ (.A1(_2156_),
    .A2(_2170_),
    .ZN(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6397_ (.A1(_2171_),
    .A2(_2176_),
    .ZN(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6398_ (.A1(_2372_),
    .A2(_2373_),
    .ZN(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6399_ (.A1(_2165_),
    .A2(_2166_),
    .B(_1957_),
    .ZN(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6400_ (.A1(_2909_),
    .A2(_2375_),
    .Z(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6401_ (.A1(_2002_),
    .A2(_1877_),
    .B(_2375_),
    .ZN(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6402_ (.A1(_2377_),
    .A2(_2378_),
    .Z(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _6403_ (.A1(_3266_),
    .A2(_1948_),
    .A3(_2163_),
    .B1(_2164_),
    .B2(_2169_),
    .ZN(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6404_ (.A1(_2347_),
    .A2(_1945_),
    .ZN(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6405_ (.A1(_2240_),
    .A2(_2198_),
    .A3(_2349_),
    .ZN(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6406_ (.A1(_2200_),
    .A2(_2381_),
    .A3(_2382_),
    .ZN(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6407_ (.A1(_2380_),
    .A2(_2383_),
    .Z(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6408_ (.A1(_2379_),
    .A2(_2384_),
    .Z(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6409_ (.A1(_2371_),
    .A2(_2374_),
    .A3(_2385_),
    .Z(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6410_ (.A1(_2152_),
    .A2(_2153_),
    .A3(_2177_),
    .ZN(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6411_ (.A1(_2152_),
    .A2(_2153_),
    .B(_2177_),
    .ZN(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6412_ (.A1(_2151_),
    .A2(_2388_),
    .B(_2389_),
    .ZN(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6413_ (.A1(_2386_),
    .A2(_2390_),
    .Z(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6414_ (.A1(_1975_),
    .A2(_1978_),
    .Z(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6415_ (.A1(_2392_),
    .A2(_2180_),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6416_ (.A1(_1935_),
    .A2(_1979_),
    .A3(_2183_),
    .B1(_2393_),
    .B2(_2182_),
    .ZN(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6417_ (.A1(_2391_),
    .A2(_2394_),
    .ZN(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6418_ (.A1(_2391_),
    .A2(_2394_),
    .Z(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6419_ (.A1(_3291_),
    .A2(_2395_),
    .A3(_2396_),
    .ZN(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6420_ (.A1(_1273_),
    .A2(_2336_),
    .A3(_2370_),
    .A4(_2397_),
    .Z(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6421_ (.I(_1269_),
    .Z(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6422_ (.A1(_2268_),
    .A2(_2301_),
    .B(_2399_),
    .C(_2400_),
    .ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6423_ (.A1(_2116_),
    .A2(_2121_),
    .ZN(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6424_ (.I(_2283_),
    .ZN(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6425_ (.A1(_2278_),
    .A2(_2402_),
    .ZN(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6426_ (.A1(_2276_),
    .A2(_2284_),
    .B(_2403_),
    .ZN(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6427_ (.A1(_2275_),
    .A2(_2401_),
    .A3(_2404_),
    .Z(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6428_ (.I(_2405_),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6429_ (.A1(_2272_),
    .A2(_2285_),
    .ZN(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6430_ (.I(_2269_),
    .ZN(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6431_ (.A1(_2409_),
    .A2(_2286_),
    .ZN(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6432_ (.A1(_2407_),
    .A2(_2410_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6433_ (.A1(_2406_),
    .A2(_2411_),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6434_ (.A1(_2407_),
    .A2(_2410_),
    .A3(_2405_),
    .ZN(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6435_ (.A1(_2412_),
    .A2(_2413_),
    .ZN(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6436_ (.A1(_2287_),
    .A2(_2292_),
    .Z(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6437_ (.A1(_2415_),
    .A2(_2300_),
    .ZN(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6438_ (.A1(_2414_),
    .A2(_2416_),
    .Z(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6439_ (.I(_1272_),
    .Z(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6440_ (.A1(_2414_),
    .A2(_2416_),
    .B(_2418_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6441_ (.A1(_2356_),
    .A2(_2360_),
    .ZN(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6442_ (.A1(_2340_),
    .A2(_2353_),
    .ZN(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6443_ (.A1(_2337_),
    .A2(_2355_),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6444_ (.A1(_2239_),
    .A2(_2241_),
    .Z(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6445_ (.I(_2351_),
    .ZN(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6446_ (.A1(_2345_),
    .A2(_2352_),
    .ZN(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6447_ (.A1(_2346_),
    .A2(_2425_),
    .B(_2426_),
    .ZN(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6448_ (.A1(_2424_),
    .A2(_2427_),
    .Z(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6449_ (.A1(_2342_),
    .A2(_2428_),
    .ZN(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6450_ (.A1(_2422_),
    .A2(_2423_),
    .B(_2429_),
    .ZN(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6451_ (.A1(_2422_),
    .A2(_2423_),
    .A3(_2429_),
    .Z(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6452_ (.A1(_2431_),
    .A2(_2432_),
    .ZN(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6453_ (.A1(_2421_),
    .A2(_2367_),
    .B(_2433_),
    .ZN(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6454_ (.A1(_2361_),
    .A2(_2366_),
    .B(_2433_),
    .C(_2421_),
    .ZN(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6455_ (.A1(_2044_),
    .A2(_2435_),
    .ZN(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6456_ (.A1(_2159_),
    .A2(_2161_),
    .Z(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6457_ (.I(_2383_),
    .ZN(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6458_ (.A1(_2379_),
    .A2(_2384_),
    .ZN(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6459_ (.A1(_2380_),
    .A2(_2438_),
    .B(_2439_),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6460_ (.A1(_2377_),
    .A2(_2437_),
    .A3(_2440_),
    .Z(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6461_ (.A1(_2374_),
    .A2(_2385_),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6462_ (.A1(_2374_),
    .A2(_2385_),
    .ZN(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6463_ (.A1(_2371_),
    .A2(_2443_),
    .B(_2444_),
    .ZN(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6464_ (.A1(_2442_),
    .A2(_2445_),
    .ZN(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6465_ (.A1(_2442_),
    .A2(_2445_),
    .Z(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6466_ (.A1(_2446_),
    .A2(_2447_),
    .ZN(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6467_ (.A1(_2386_),
    .A2(_2390_),
    .ZN(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6468_ (.A1(_2391_),
    .A2(_2394_),
    .B(_2449_),
    .ZN(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6469_ (.A1(_2448_),
    .A2(_2450_),
    .Z(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6470_ (.I(_2145_),
    .Z(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6471_ (.A1(_2434_),
    .A2(_2436_),
    .B1(_2451_),
    .B2(_2453_),
    .ZN(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6472_ (.A1(_2305_),
    .A2(_2315_),
    .ZN(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6473_ (.I(_2455_),
    .ZN(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6474_ (.A1(_2302_),
    .A2(_2316_),
    .Z(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6475_ (.A1(_2199_),
    .A2(_2202_),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6476_ (.I(_2313_),
    .ZN(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6477_ (.A1(_2311_),
    .A2(_2459_),
    .ZN(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6478_ (.A1(_2309_),
    .A2(_2314_),
    .B(_2460_),
    .ZN(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6479_ (.A1(_2308_),
    .A2(_2458_),
    .A3(_2461_),
    .Z(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6480_ (.I(_2462_),
    .ZN(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6481_ (.A1(_2456_),
    .A2(_2457_),
    .B(_2464_),
    .ZN(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6482_ (.A1(_2456_),
    .A2(_2457_),
    .A3(_2464_),
    .Z(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6483_ (.A1(_2465_),
    .A2(_2466_),
    .ZN(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6484_ (.A1(_2317_),
    .A2(_2322_),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6485_ (.A1(_2323_),
    .A2(_2333_),
    .B(_2468_),
    .ZN(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6486_ (.A1(_2467_),
    .A2(_2469_),
    .Z(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6487_ (.A1(_1271_),
    .A2(_2470_),
    .B(_3296_),
    .ZN(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6488_ (.A1(_2417_),
    .A2(_2420_),
    .B1(_2454_),
    .B2(_2471_),
    .C(_2266_),
    .ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6489_ (.A1(_2415_),
    .A2(_2412_),
    .ZN(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6490_ (.A1(_2401_),
    .A2(_2404_),
    .ZN(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6491_ (.A1(_2401_),
    .A2(_2404_),
    .ZN(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6492_ (.A1(_2275_),
    .A2(_2474_),
    .B(_2475_),
    .C(_2264_),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6493_ (.A1(_2300_),
    .A2(_2414_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6494_ (.A1(_2413_),
    .A2(_2472_),
    .B(_2476_),
    .C(_2477_),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6495_ (.A1(_2437_),
    .A2(_2440_),
    .ZN(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6496_ (.A1(_2437_),
    .A2(_2440_),
    .ZN(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6497_ (.A1(_2377_),
    .A2(_2479_),
    .B(_2480_),
    .ZN(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6498_ (.A1(_2446_),
    .A2(_2481_),
    .ZN(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6499_ (.A1(_2449_),
    .A2(_2447_),
    .B(_2482_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6500_ (.A1(_2395_),
    .A2(_2448_),
    .B(_2483_),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6501_ (.A1(_2458_),
    .A2(_2461_),
    .ZN(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6502_ (.A1(_2458_),
    .A2(_2461_),
    .ZN(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6503_ (.A1(_2308_),
    .A2(_2486_),
    .B(_2465_),
    .C(_2487_),
    .ZN(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6504_ (.A1(_2468_),
    .A2(_2466_),
    .B(_2488_),
    .ZN(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6505_ (.A1(_2334_),
    .A2(_2467_),
    .B(_2489_),
    .ZN(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6506_ (.I(_1924_),
    .Z(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6507_ (.A1(_2361_),
    .A2(_2366_),
    .A3(_2433_),
    .ZN(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6508_ (.I(_2432_),
    .ZN(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6509_ (.A1(_2342_),
    .A2(_2428_),
    .ZN(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6510_ (.A1(_2424_),
    .A2(_2427_),
    .B(_2494_),
    .C(_1923_),
    .ZN(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6511_ (.A1(_2421_),
    .A2(_2493_),
    .B(_2496_),
    .C(_2431_),
    .ZN(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6512_ (.A1(_2492_),
    .A2(_2497_),
    .B(_2225_),
    .ZN(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6513_ (.A1(_2147_),
    .A2(_2485_),
    .B1(_2490_),
    .B2(_2491_),
    .C(_2498_),
    .ZN(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6514_ (.A1(_2400_),
    .A2(_2478_),
    .A3(_2499_),
    .ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6515_ (.I(_2264_),
    .Z(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6516_ (.A1(_3186_),
    .A2(_2453_),
    .ZN(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6517_ (.A1(_3103_),
    .A2(_3185_),
    .B(_2501_),
    .ZN(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6518_ (.A1(_0490_),
    .A2(_0407_),
    .B1(_0472_),
    .B2(_0491_),
    .ZN(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6519_ (.A1(_1069_),
    .A2(_1157_),
    .ZN(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6520_ (.A1(_2368_),
    .A2(_2504_),
    .ZN(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6521_ (.A1(_0492_),
    .A2(_2226_),
    .A3(_2503_),
    .B1(_2506_),
    .B2(_1159_),
    .ZN(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6522_ (.A1(_1731_),
    .A2(_0490_),
    .B1(_1772_),
    .B2(_0491_),
    .ZN(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6523_ (.A1(_1788_),
    .A2(_2508_),
    .B(_2101_),
    .ZN(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6524_ (.A1(_2500_),
    .A2(_2502_),
    .A3(_2507_),
    .B(_2509_),
    .ZN(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6525_ (.A1(_2400_),
    .A2(_2510_),
    .ZN(net17));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6526_ (.A1(_1718_),
    .A2(_1787_),
    .A3(_1788_),
    .Z(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6527_ (.A1(_3076_),
    .A2(_3187_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6528_ (.A1(_3188_),
    .A2(_3291_),
    .A3(_2512_),
    .ZN(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6529_ (.A1(_1044_),
    .A2(_1161_),
    .B(_2043_),
    .ZN(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6530_ (.A1(_0388_),
    .A2(_0489_),
    .A3(_0492_),
    .ZN(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6531_ (.A1(_1162_),
    .A2(_2514_),
    .B1(_2516_),
    .B2(_1925_),
    .ZN(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6532_ (.A1(_2418_),
    .A2(_2513_),
    .A3(_2517_),
    .Z(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6533_ (.A1(_2268_),
    .A2(_2511_),
    .B(_2518_),
    .C(_2400_),
    .ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6534_ (.A1(_0495_),
    .A2(_0496_),
    .Z(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6535_ (.A1(_0497_),
    .A2(_2491_),
    .A3(_2519_),
    .ZN(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6536_ (.A1(_1163_),
    .A2(_1164_),
    .B(_2044_),
    .ZN(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6537_ (.A1(_3189_),
    .A2(_3190_),
    .B(_2145_),
    .ZN(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6538_ (.A1(_3191_),
    .A2(_2522_),
    .B(_1273_),
    .ZN(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6539_ (.A1(_1165_),
    .A2(_2521_),
    .B(_2523_),
    .ZN(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6540_ (.A1(_1786_),
    .A2(_1791_),
    .ZN(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6541_ (.A1(_2520_),
    .A2(_2524_),
    .B1(_2526_),
    .B2(_2103_),
    .C(_2266_),
    .ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6542_ (.A1(_1784_),
    .A2(_1792_),
    .ZN(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6543_ (.A1(_0487_),
    .A2(_0497_),
    .B(_2226_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6544_ (.A1(_3180_),
    .A2(_3191_),
    .Z(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6545_ (.A1(_3180_),
    .A2(_3191_),
    .B(_2145_),
    .ZN(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6546_ (.A1(_1153_),
    .A2(_1165_),
    .ZN(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6547_ (.A1(_1166_),
    .A2(_2368_),
    .A3(_2531_),
    .ZN(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6548_ (.A1(_2529_),
    .A2(_2530_),
    .B(_2532_),
    .C(_1273_),
    .ZN(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6549_ (.A1(_0498_),
    .A2(_2528_),
    .B(_2533_),
    .ZN(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6550_ (.A1(_2268_),
    .A2(_2527_),
    .B(_2534_),
    .C(_1270_),
    .ZN(net27));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6551_ (.A1(_0470_),
    .A2(_0502_),
    .Z(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6552_ (.A1(_0498_),
    .A2(_2536_),
    .ZN(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6553_ (.A1(_0499_),
    .A2(_2491_),
    .A3(_2537_),
    .ZN(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6554_ (.A1(_3166_),
    .A2(_3195_),
    .Z(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6555_ (.A1(_2529_),
    .A2(_2539_),
    .ZN(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6556_ (.A1(_1981_),
    .A2(_2540_),
    .ZN(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6557_ (.A1(_1137_),
    .A2(_1151_),
    .ZN(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6558_ (.A1(_1166_),
    .A2(_2542_),
    .B(_2044_),
    .C(_1167_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6559_ (.A1(_3193_),
    .A2(_2541_),
    .B(_2543_),
    .C(_2500_),
    .ZN(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6560_ (.I(_1267_),
    .Z(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6561_ (.A1(_1749_),
    .A2(_1759_),
    .Z(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6562_ (.A1(_1766_),
    .A2(_1780_),
    .ZN(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6563_ (.A1(_1784_),
    .A2(_1792_),
    .ZN(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6564_ (.A1(_2547_),
    .A2(_2548_),
    .A3(_2549_),
    .ZN(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6565_ (.A1(_1793_),
    .A2(_1781_),
    .A3(_2550_),
    .B(_0696_),
    .ZN(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6566_ (.A1(_2546_),
    .A2(_2551_),
    .ZN(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6567_ (.A1(_2538_),
    .A2(_2544_),
    .B(_2552_),
    .ZN(net28));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6568_ (.A1(_3193_),
    .A2(_3198_),
    .ZN(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6569_ (.A1(_3199_),
    .A2(_2147_),
    .A3(_2553_),
    .ZN(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6570_ (.A1(_0499_),
    .A2(_0505_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6571_ (.A1(_0506_),
    .A2(_2226_),
    .ZN(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6572_ (.A1(_1167_),
    .A2(_1171_),
    .B(_2368_),
    .ZN(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6573_ (.A1(_1172_),
    .A2(_2558_),
    .B(_2418_),
    .ZN(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6574_ (.A1(_2556_),
    .A2(_2557_),
    .B(_2559_),
    .ZN(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6575_ (.A1(_1793_),
    .A2(_1783_),
    .Z(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6576_ (.A1(_1274_),
    .A2(_2561_),
    .B(_2546_),
    .ZN(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6577_ (.A1(_2554_),
    .A2(_2560_),
    .B(_2562_),
    .ZN(net29));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6578_ (.A1(_1794_),
    .A2(_1795_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6579_ (.A1(_0506_),
    .A2(_0507_),
    .A3(_0510_),
    .ZN(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6580_ (.A1(_0506_),
    .A2(_0507_),
    .B(_0510_),
    .ZN(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6581_ (.A1(_2566_),
    .A2(_1925_),
    .ZN(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6582_ (.A1(_2564_),
    .A2(_2567_),
    .B(_2418_),
    .ZN(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6583_ (.A1(_3201_),
    .A2(_3204_),
    .Z(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6584_ (.A1(_3201_),
    .A2(_3204_),
    .ZN(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6585_ (.A1(_2569_),
    .A2(_2453_),
    .A3(_2570_),
    .ZN(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6586_ (.A1(_1173_),
    .A2(_1176_),
    .Z(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6587_ (.A1(_1173_),
    .A2(_1176_),
    .ZN(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6588_ (.A1(_2572_),
    .A2(_0585_),
    .A3(_2573_),
    .ZN(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6589_ (.A1(_2571_),
    .A2(_2574_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6590_ (.A1(_2568_),
    .A2(_2575_),
    .B(_2546_),
    .ZN(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6591_ (.A1(_2268_),
    .A2(_2563_),
    .B(_2577_),
    .ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6592_ (.A1(_1747_),
    .A2(_1799_),
    .ZN(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6593_ (.A1(_0508_),
    .A2(_0509_),
    .ZN(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6594_ (.A1(_2579_),
    .A2(_2566_),
    .ZN(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6595_ (.A1(_0452_),
    .A2(_0459_),
    .A3(_2580_),
    .Z(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6596_ (.A1(_3147_),
    .A2(_3209_),
    .Z(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6597_ (.A1(_3206_),
    .A2(_2569_),
    .B(_2582_),
    .ZN(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6598_ (.A1(_3206_),
    .A2(_2569_),
    .A3(_2582_),
    .Z(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6599_ (.A1(_1178_),
    .A2(_2572_),
    .ZN(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6600_ (.A1(_1115_),
    .A2(_1182_),
    .A3(_2585_),
    .Z(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6601_ (.A1(_1981_),
    .A2(_2583_),
    .A3(_2584_),
    .B1(_2587_),
    .B2(_2225_),
    .ZN(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6602_ (.A1(_3296_),
    .A2(_2581_),
    .B(_2588_),
    .C(_2101_),
    .ZN(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6603_ (.A1(_2103_),
    .A2(_2578_),
    .B(_2589_),
    .C(_1270_),
    .ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6604_ (.A1(_1714_),
    .A2(_1801_),
    .Z(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6605_ (.A1(_1714_),
    .A2(_1801_),
    .ZN(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6606_ (.A1(_2590_),
    .A2(_2591_),
    .ZN(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6607_ (.A1(_3210_),
    .A2(_3214_),
    .Z(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6608_ (.A1(_3210_),
    .A2(_3214_),
    .ZN(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6609_ (.A1(_2593_),
    .A2(_2453_),
    .A3(_2594_),
    .ZN(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6610_ (.A1(_1183_),
    .A2(_1187_),
    .Z(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6611_ (.A1(_1183_),
    .A2(_1187_),
    .B(_2043_),
    .ZN(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6612_ (.A1(_0514_),
    .A2(_0519_),
    .Z(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6613_ (.A1(_2597_),
    .A2(_2598_),
    .B1(_2599_),
    .B2(_2491_),
    .C(_2264_),
    .ZN(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6614_ (.A1(_2103_),
    .A2(_2592_),
    .B1(_2595_),
    .B2(_2600_),
    .C(_2266_),
    .ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6615_ (.A1(_3211_),
    .A2(_3213_),
    .B(_2593_),
    .ZN(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6616_ (.A1(_3070_),
    .A2(_2601_),
    .ZN(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6617_ (.A1(_2147_),
    .A2(_2602_),
    .B(_2500_),
    .ZN(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6618_ (.A1(_0515_),
    .A2(_0518_),
    .ZN(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6619_ (.A1(_0514_),
    .A2(_0519_),
    .ZN(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6620_ (.A1(_2604_),
    .A2(_2605_),
    .ZN(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6621_ (.A1(_0383_),
    .A2(_2607_),
    .Z(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6622_ (.A1(_1184_),
    .A2(_1186_),
    .B(_2597_),
    .ZN(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6623_ (.A1(_1036_),
    .A2(_2609_),
    .Z(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6624_ (.A1(_2225_),
    .A2(_2610_),
    .ZN(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6625_ (.A1(_3296_),
    .A2(_2608_),
    .B(_2611_),
    .ZN(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6626_ (.A1(_1803_),
    .A2(_2590_),
    .ZN(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6627_ (.A1(_1659_),
    .A2(_1660_),
    .A3(_2613_),
    .Z(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6628_ (.A1(_1274_),
    .A2(_2614_),
    .B(_2546_),
    .ZN(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6629_ (.A1(_2603_),
    .A2(_2612_),
    .B(_2615_),
    .ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6630_ (.A1(_1661_),
    .A2(_1804_),
    .B(_1586_),
    .ZN(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6631_ (.A1(_1805_),
    .A2(_2617_),
    .Z(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6632_ (.A1(_1194_),
    .A2(_1188_),
    .A3(_1193_),
    .Z(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6633_ (.A1(_1195_),
    .A2(_0585_),
    .A3(_2619_),
    .ZN(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6634_ (.A1(_0304_),
    .A2(_0525_),
    .B(_1924_),
    .ZN(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6635_ (.A1(_0304_),
    .A2(_0525_),
    .B(_2621_),
    .ZN(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6636_ (.A1(_3220_),
    .A2(_3215_),
    .A3(_3218_),
    .ZN(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6637_ (.A1(_3221_),
    .A2(_3291_),
    .ZN(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6638_ (.A1(_2623_),
    .A2(_2624_),
    .ZN(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6639_ (.A1(_2101_),
    .A2(_2622_),
    .A3(_2625_),
    .ZN(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6640_ (.A1(_2500_),
    .A2(_2618_),
    .B1(_2620_),
    .B2(_2626_),
    .C(_1269_),
    .ZN(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6641_ (.I(net3),
    .Z(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6642_ (.A1(net2),
    .A2(net12),
    .ZN(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6643_ (.A1(net14),
    .A2(net13),
    .ZN(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6644_ (.A1(_2629_),
    .A2(_2630_),
    .Z(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6645_ (.I(_2631_),
    .Z(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6646_ (.I0(_0490_),
    .I1(_2628_),
    .S(_2632_),
    .Z(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6647_ (.I(_2633_),
    .Z(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6648_ (.I(net4),
    .Z(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6649_ (.I0(_0350_),
    .I1(_2634_),
    .S(_2632_),
    .Z(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6650_ (.I(_2635_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6651_ (.I(net5),
    .Z(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6652_ (.I(_2631_),
    .Z(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6653_ (.I0(_0547_),
    .I1(_2637_),
    .S(_2638_),
    .Z(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6654_ (.I(_2639_),
    .Z(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6655_ (.I(net6),
    .Z(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6656_ (.I0(_0548_),
    .I1(_2640_),
    .S(_2638_),
    .Z(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6657_ (.I(_2641_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6658_ (.I(net7),
    .Z(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6659_ (.I0(_1437_),
    .I1(_2642_),
    .S(_2638_),
    .Z(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6660_ (.I(_2643_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6661_ (.I(net8),
    .Z(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6662_ (.I0(_2118_),
    .I1(_2645_),
    .S(_2638_),
    .Z(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6663_ (.I(_2646_),
    .Z(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6664_ (.I(net9),
    .Z(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6665_ (.I0(_2119_),
    .I1(_2647_),
    .S(_2631_),
    .Z(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6666_ (.I(_2648_),
    .Z(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6667_ (.I(net10),
    .Z(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6668_ (.A1(_2649_),
    .A2(_2632_),
    .ZN(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6669_ (.A1(_2279_),
    .A2(_2632_),
    .B(_2650_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6670_ (.I(net3),
    .Z(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6671_ (.I(net12),
    .ZN(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6672_ (.A1(net2),
    .A2(_2653_),
    .ZN(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6673_ (.A1(_2630_),
    .A2(_2654_),
    .ZN(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6674_ (.I(_2655_),
    .Z(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6675_ (.I0(_2652_),
    .I1(_0491_),
    .S(_2656_),
    .Z(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6676_ (.I(_2657_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6677_ (.I(net4),
    .Z(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6678_ (.I0(_2658_),
    .I1(_0473_),
    .S(_2656_),
    .Z(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6679_ (.I(_2659_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6680_ (.I(net5),
    .Z(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6681_ (.I0(_2661_),
    .I1(_0191_),
    .S(_2656_),
    .Z(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6682_ (.I(_2662_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6683_ (.I(net6),
    .Z(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6684_ (.I0(_2663_),
    .I1(_0530_),
    .S(_2656_),
    .Z(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6685_ (.I(_2664_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6686_ (.I(net7),
    .Z(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6687_ (.I(_2655_),
    .Z(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6688_ (.I0(_2665_),
    .I1(_1817_),
    .S(_2666_),
    .Z(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6689_ (.I(_2667_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6690_ (.I(net8),
    .Z(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6691_ (.I0(_2669_),
    .I1(_1612_),
    .S(_2666_),
    .Z(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6692_ (.I(_2670_),
    .Z(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6693_ (.I(net9),
    .Z(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6694_ (.I0(_2671_),
    .I1(_2131_),
    .S(_2666_),
    .Z(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6695_ (.I(_2672_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6696_ (.I(net10),
    .Z(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6697_ (.I0(_2673_),
    .I1(_2058_),
    .S(_2666_),
    .Z(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6698_ (.I(_2674_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6699_ (.I(net13),
    .ZN(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6700_ (.A1(net14),
    .A2(_2675_),
    .ZN(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6701_ (.A1(_2629_),
    .A2(_2677_),
    .ZN(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6702_ (.I(_2678_),
    .Z(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6703_ (.I0(_2652_),
    .I1(_3102_),
    .S(_2679_),
    .Z(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6704_ (.I(_2680_),
    .Z(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6705_ (.I0(_2658_),
    .I1(_2933_),
    .S(_2679_),
    .Z(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6706_ (.I(_2681_),
    .Z(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6707_ (.I(_2678_),
    .Z(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6708_ (.I0(_2661_),
    .I1(_3246_),
    .S(_2682_),
    .Z(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6709_ (.I(_2683_),
    .Z(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6710_ (.I0(_2663_),
    .I1(_3247_),
    .S(_2682_),
    .Z(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6711_ (.I(_2685_),
    .Z(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6712_ (.I0(_2665_),
    .I1(_3272_),
    .S(_2682_),
    .Z(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6713_ (.I(_2686_),
    .Z(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6714_ (.I0(_2669_),
    .I1(_2160_),
    .S(_2682_),
    .Z(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6715_ (.I(_2687_),
    .Z(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6716_ (.I0(_2671_),
    .I1(_2240_),
    .S(_2678_),
    .Z(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6717_ (.I(_2688_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6718_ (.A1(_2649_),
    .A2(_2679_),
    .ZN(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6719_ (.A1(_2347_),
    .A2(_2679_),
    .B(_2689_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6720_ (.A1(_2654_),
    .A2(_2677_),
    .ZN(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6721_ (.I(_2691_),
    .Z(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6722_ (.I0(_2652_),
    .I1(_3025_),
    .S(_2692_),
    .Z(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6723_ (.I(_2693_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6724_ (.I0(_2658_),
    .I1(_1829_),
    .S(_2692_),
    .Z(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6725_ (.I(_2694_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6726_ (.I0(_2661_),
    .I1(_2910_),
    .S(_2692_),
    .Z(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6727_ (.I(_2695_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6728_ (.I0(_2663_),
    .I1(_3225_),
    .S(_2692_),
    .Z(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6729_ (.I(_2696_),
    .Z(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6730_ (.I(_2691_),
    .Z(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6731_ (.I0(_2665_),
    .I1(_1208_),
    .S(_2698_),
    .Z(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6732_ (.I(_2699_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6733_ (.I0(_2669_),
    .I1(_0979_),
    .S(_2698_),
    .Z(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6734_ (.I(_2700_),
    .Z(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6735_ (.I0(_2671_),
    .I1(_2003_),
    .S(_2698_),
    .Z(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6736_ (.I(_2701_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6737_ (.I0(_2673_),
    .I1(_2002_),
    .S(_2698_),
    .Z(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6738_ (.I(_2702_),
    .Z(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6739_ (.A1(net14),
    .A2(_2675_),
    .Z(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6740_ (.A1(_2629_),
    .A2(_2703_),
    .ZN(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6741_ (.I(_2705_),
    .Z(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6742_ (.I0(_2652_),
    .I1(_1731_),
    .S(_2706_),
    .Z(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6743_ (.I(_2707_),
    .Z(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6744_ (.I0(_2658_),
    .I1(_1140_),
    .S(_2706_),
    .Z(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6745_ (.I(_2708_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6746_ (.I0(_2661_),
    .I1(_1007_),
    .S(_2706_),
    .Z(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6747_ (.I(_2709_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6748_ (.I0(_2663_),
    .I1(_0998_),
    .S(_2706_),
    .Z(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6749_ (.I(_2710_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6750_ (.I(_2705_),
    .Z(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6751_ (.I0(_2665_),
    .I1(_1000_),
    .S(_2712_),
    .Z(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6752_ (.I(_2713_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6753_ (.I0(_2669_),
    .I1(_1241_),
    .S(_2712_),
    .Z(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6754_ (.I(_2714_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6755_ (.I0(_2671_),
    .I1(_2117_),
    .S(_2712_),
    .Z(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6756_ (.I(_2715_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6757_ (.I0(_2673_),
    .I1(_2120_),
    .S(_2712_),
    .Z(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6758_ (.I(_2716_),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6759_ (.A1(_2654_),
    .A2(_2703_),
    .ZN(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6760_ (.I(_2717_),
    .Z(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6761_ (.I0(_2628_),
    .I1(_0407_),
    .S(_2719_),
    .Z(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6762_ (.I(_2720_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6763_ (.I0(_2634_),
    .I1(_3169_),
    .S(_2719_),
    .Z(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6764_ (.I(_2721_),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6765_ (.I0(_2637_),
    .I1(_3098_),
    .S(_2719_),
    .Z(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6766_ (.I(_2722_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6767_ (.I0(_2640_),
    .I1(_3032_),
    .S(_2719_),
    .Z(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6768_ (.I(_2723_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6769_ (.I(_2717_),
    .Z(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6770_ (.I0(_2642_),
    .I1(_3034_),
    .S(_2724_),
    .Z(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6771_ (.I(_2726_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6772_ (.I0(_2645_),
    .I1(_3262_),
    .S(_2724_),
    .Z(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6773_ (.I(_2727_),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6774_ (.I0(_2647_),
    .I1(_2198_),
    .S(_2724_),
    .Z(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6775_ (.I(_2728_),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6776_ (.I0(_2673_),
    .I1(_2200_),
    .S(_2724_),
    .Z(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6777_ (.I(_2729_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6778_ (.A1(net14),
    .A2(net13),
    .ZN(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6779_ (.A1(_1267_),
    .A2(net12),
    .A3(_2730_),
    .ZN(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6780_ (.I(_2731_),
    .Z(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6781_ (.I0(_1772_),
    .I1(_2628_),
    .S(_2733_),
    .Z(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6782_ (.I(_2734_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6783_ (.I0(_1043_),
    .I1(_2634_),
    .S(_2733_),
    .Z(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6784_ (.I(_2735_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6785_ (.I0(_1039_),
    .I1(_2637_),
    .S(_2733_),
    .Z(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6786_ (.I(_2736_),
    .Z(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6787_ (.I0(_0830_),
    .I1(_2640_),
    .S(_2733_),
    .Z(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6788_ (.I(_2737_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6789_ (.I(_2731_),
    .Z(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6790_ (.I0(_1596_),
    .I1(_2642_),
    .S(_2738_),
    .Z(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6791_ (.I(_2740_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6792_ (.I0(_1595_),
    .I1(_2645_),
    .S(_2738_),
    .Z(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6793_ (.I(_2741_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6794_ (.I0(_2005_),
    .I1(_2647_),
    .S(_2738_),
    .Z(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6795_ (.I(_2742_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6796_ (.I0(_1811_),
    .I1(_2649_),
    .S(_2738_),
    .Z(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6797_ (.I(_2743_),
    .Z(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6798_ (.A1(_1267_),
    .A2(_2653_),
    .A3(_2730_),
    .ZN(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6799_ (.I(_2744_),
    .Z(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6800_ (.I0(_0472_),
    .I1(_2628_),
    .S(_2745_),
    .Z(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6801_ (.I(_2747_),
    .Z(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6802_ (.I0(_3075_),
    .I1(_2634_),
    .S(_2745_),
    .Z(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6803_ (.I(_2748_),
    .Z(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6804_ (.I0(_3174_),
    .I1(_2637_),
    .S(_2745_),
    .Z(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6805_ (.I(_2749_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6806_ (.I0(_2940_),
    .I1(_2640_),
    .S(_2745_),
    .Z(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6807_ (.I(_2750_),
    .Z(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6808_ (.I(_2744_),
    .Z(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6809_ (.I0(_0319_),
    .I1(_2642_),
    .S(_2751_),
    .Z(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6810_ (.I(_2752_),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6811_ (.I0(_0317_),
    .I1(_2645_),
    .S(_2751_),
    .Z(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6812_ (.I(_2754_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6813_ (.I0(_1898_),
    .I1(_2647_),
    .S(_2751_),
    .Z(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6814_ (.I(_2755_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6815_ (.I0(_1877_),
    .I1(_2649_),
    .S(_2751_),
    .Z(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6816_ (.I(_2756_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6817_ (.D(_0000_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6818_ (.D(_0001_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6819_ (.D(_0002_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6820_ (.D(_0003_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6821_ (.D(_0004_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6822_ (.D(_0005_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6823_ (.D(_0006_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6824_ (.D(_0007_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6825_ (.D(_0008_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6826_ (.D(_0009_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6827_ (.D(_0010_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6828_ (.D(_0011_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6829_ (.D(_0012_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6830_ (.D(_0013_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6831_ (.D(_0014_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6832_ (.D(_0015_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6833_ (.D(_0016_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6834_ (.D(_0017_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6835_ (.D(_0018_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6836_ (.D(_0019_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6837_ (.D(_0020_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6838_ (.D(_0021_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6839_ (.D(_0022_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6840_ (.D(_0023_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6841_ (.D(_0024_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6842_ (.D(_0025_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6843_ (.D(_0026_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6844_ (.D(_0027_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6845_ (.D(_0028_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6846_ (.D(_0029_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6847_ (.D(_0030_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6848_ (.D(_0031_),
    .RN(net11),
    .CLK(net1),
    .Q(\A[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6849_ (.D(_0032_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6850_ (.D(_0033_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6851_ (.D(_0034_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6852_ (.D(_0035_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6853_ (.D(_0036_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6854_ (.D(_0037_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6855_ (.D(_0038_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6856_ (.D(_0039_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6857_ (.D(_0040_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6858_ (.D(_0041_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6859_ (.D(_0042_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6860_ (.D(_0043_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6861_ (.D(_0044_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6862_ (.D(_0045_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6863_ (.D(_0046_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6864_ (.D(_0047_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6865_ (.D(_0048_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6866_ (.D(_0049_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6867_ (.D(_0050_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6868_ (.D(_0051_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6869_ (.D(_0052_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6870_ (.D(_0053_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6871_ (.D(_0054_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6872_ (.D(_0055_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6873_ (.D(_0056_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6874_ (.D(_0057_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6875_ (.D(_0058_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6876_ (.D(_0059_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6877_ (.D(_0060_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6878_ (.D(_0061_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6879_ (.D(_0062_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _6880_ (.D(_0063_),
    .RN(net11),
    .CLK(net1),
    .Q(\B[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 input1 (.I(clk),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(execute),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(input_val[0]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(input_val[1]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(input_val[2]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(input_val[3]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(input_val[4]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(input_val[5]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(input_val[6]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(input_val[7]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_20 input11 (.I(reset),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(sel_in[0]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(sel_in[1]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input14 (.I(sel_in[2]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(sel_out[0]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(sel_out[1]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output17 (.I(net17),
    .Z(result[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output18 (.I(net18),
    .Z(result[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output19 (.I(net19),
    .Z(result[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output20 (.I(net20),
    .Z(result[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output21 (.I(net21),
    .Z(result[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output22 (.I(net22),
    .Z(result[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output23 (.I(net23),
    .Z(result[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output24 (.I(net24),
    .Z(result[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output25 (.I(net25),
    .Z(result[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output26 (.I(net26),
    .Z(result[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output27 (.I(net27),
    .Z(result[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output28 (.I(net28),
    .Z(result[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output29 (.I(net29),
    .Z(result[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output30 (.I(net30),
    .Z(result[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output31 (.I(net31),
    .Z(result[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output32 (.I(net32),
    .Z(result[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output33 (.I(net33),
    .Z(result[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4503__I (.I(\A[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__A2 (.I(\A[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__A3 (.I(\A[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4168__I (.I(\A[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A1 (.I(\A[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__B1 (.I(\A[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__A4 (.I(\A[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__I (.I(\A[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A2 (.I(\A[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__A2 (.I(\A[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__I (.I(\A[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__I (.I(\A[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__A1 (.I(\A[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A1 (.I(\A[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4185__I (.I(\A[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__A1 (.I(\A[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A1 (.I(\A[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4190__I (.I(\A[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__I (.I(\A[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__I (.I(\A[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__A1 (.I(\A[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__I (.I(\A[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__A1 (.I(\A[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A3 (.I(\A[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__A2 (.I(\A[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__A3 (.I(\A[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3452__I (.I(\A[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3566__I (.I(\A[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3528__I (.I(\A[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3516__I (.I(\A[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A1 (.I(\A[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3732__I (.I(\A[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A1 (.I(\A[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3593__I (.I(\A[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3470__I (.I(\A[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3434__I (.I(\A[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3475__I (.I(\A[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3461__I (.I(\A[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__A1 (.I(\A[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__I (.I(\A[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__I (.I(\A[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__A2 (.I(\B[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__I (.I(\B[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__I (.I(\B[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__A2 (.I(\B[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__I (.I(\B[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__I (.I(\B[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A2 (.I(\B[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__I (.I(\B[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__I (.I(\B[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3536__I (.I(\B[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3530__I (.I(\B[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3518__I (.I(\B[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A2 (.I(\B[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A2 (.I(\B[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3581__I (.I(\B[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3444__I (.I(\B[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A2 (.I(\B[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__A2 (.I(\B[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3548__I (.I(\B[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3447__I (.I(\B[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A2 (.I(\B[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__I (.I(\B[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__A2 (.I(\B[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__I (.I(\B[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__I (.I(\B[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__A2 (.I(\B[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__I (.I(\B[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__I (.I(\B[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__I (.I(\B[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__A2 (.I(\B[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3465__I (.I(\B[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A2 (.I(\B[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__A2 (.I(\B[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3484__I (.I(\B[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3407__I (.I(\B[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__A1 (.I(\B[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3486__I (.I(\B[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3409__I (.I(\B[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__D (.I(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__D (.I(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__D (.I(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__D (.I(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__D (.I(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A1 (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A2 (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__I (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A2 (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__A2 (.I(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__B1 (.I(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__A2 (.I(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__I (.I(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A2 (.I(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__I (.I(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A2 (.I(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__A2 (.I(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__A1 (.I(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A1 (.I(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__A1 (.I(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4249__I (.I(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A1 (.I(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A1 (.I(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A1 (.I(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__A1 (.I(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__A1 (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__A2 (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__I (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A1 (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A1 (.I(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A1 (.I(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__A2 (.I(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4256__I (.I(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__A1 (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A1 (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A1 (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A1 (.I(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__A2 (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4262__A2 (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__A2 (.I(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__A1 (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A1 (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A1 (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A2 (.I(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__A2 (.I(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A2 (.I(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__A1 (.I(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4301__A1 (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__A1 (.I(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4322__A1 (.I(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4272__B (.I(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A1 (.I(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A1 (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A1 (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A2 (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A1 (.I(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A1 (.I(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A1 (.I(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__A1 (.I(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A1 (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__A1 (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A1 (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__A1 (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A2 (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A4 (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A1 (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4288__I (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__A1 (.I(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__B1 (.I(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__B2 (.I(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A2 (.I(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A2 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A2 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A4 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__A2 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A2 (.I(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A2 (.I(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4294__A3 (.I(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__A2 (.I(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A2 (.I(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A2 (.I(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A1 (.I(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__A1 (.I(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__A2 (.I(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A3 (.I(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__A2 (.I(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5484__A2 (.I(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A1 (.I(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A2 (.I(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A1 (.I(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__I (.I(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__B2 (.I(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A1 (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__A1 (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A1 (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A1 (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A2 (.I(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__A2 (.I(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__A3 (.I(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A1 (.I(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__A1 (.I(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__A2 (.I(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__B1 (.I(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__A1 (.I(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__I (.I(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__B2 (.I(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A1 (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4374__A1 (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__A1 (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A3 (.I(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__I (.I(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A3 (.I(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__A2 (.I(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__A2 (.I(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__A1 (.I(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A4 (.I(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__A2 (.I(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__A1 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__A1 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__I (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A1 (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A2 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__B2 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__I (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__B2 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A2 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__A2 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__A2 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__A2 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__A2 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__A2 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A2 (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__A2 (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__A1 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__A1 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__A2 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__A2 (.I(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A2 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__A1 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__A2 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__I (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A2 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A2 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A2 (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4367__I (.I(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__I1 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A2 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__A2 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A2 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__B (.I(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__A1 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A1 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A1 (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__A1 (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__A1 (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__A1 (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__B (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A1 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__A1 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A1 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__A1 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A2 (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__A1 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4401__A1 (.I(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__A2 (.I(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__A2 (.I(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__I (.I(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A2 (.I(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A1 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__A1 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__A1 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__I (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A1 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A1 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A1 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__A2 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__A3 (.I(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__A2 (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__A2 (.I(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__A2 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A2 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__A2 (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A2 (.I(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__A2 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A2 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__B1 (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__I (.I(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__B1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__A2 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__B1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__I (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__A2 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__I (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A2 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__A2 (.I(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A1 (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A1 (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A1 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__A1 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4447__A2 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__A1 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A2 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A2 (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A1 (.I(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A2 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4458__I (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__A1 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4526__I (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__A2 (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A2 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A1 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__A1 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__A1 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__I (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__I (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__A1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__A1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A2 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A1 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A1 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__A2 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__A3 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__A2 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A2 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__A1 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6634__A1 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__A1 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A1 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A2 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__I (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A1 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__A2 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4563__I (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__I (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A2 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__A1 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__A3 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A1 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A3 (.I(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A1 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__I (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6811__I0 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A2 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A2 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__A1 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A2 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__I (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__A2 (.I(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6809__I0 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A2 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A2 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__B2 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__I (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__A2 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__I (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__A1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__A1 (.I(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__A1 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__A2 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__I (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__B2 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__A1 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__I (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A1 (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__A3 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__A3 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__A4 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4510__A2 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A4 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__A2 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__A1 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__A2 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__I0 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__A3 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A3 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__A1 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__A2 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__I (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__B2 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A3 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__B1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__A2 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A4 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__B2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__B1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A2 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A2 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A2 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A2 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__A2 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4545__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__A2 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__A3 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__A1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__I (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__B2 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__A2 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A1 (.I(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A1 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A2 (.I(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__A2 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__I (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A1 (.I(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__A1 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A2 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__A2 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__A2 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6761__I1 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A3 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__I (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A2 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__A2 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A2 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__A1 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A1 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A2 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__A2 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A1 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__A2 (.I(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__A2 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A2 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__A3 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__A1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__I (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__A2 (.I(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A2 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A2 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__A3 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A2 (.I(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A1 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A1 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A2 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A2 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A3 (.I(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A3 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A2 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__A2 (.I(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A2 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A2 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6595__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__B (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A1 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A3 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__A2 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A2 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4642__A2 (.I(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__I0 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__B1 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A4 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A1 (.I(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__I1 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A2 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A2 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A2 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__I (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__A1 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A3 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A4 (.I(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6646__I0 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__A1 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A1 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__I1 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__B2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__B2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__A3 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A2 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__B1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6619__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__A2 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__A2 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__B3 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__A2 (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A2 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__A2 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__A2 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6634__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__B (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__I1 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A2 (.I(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A1 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__B1 (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A4 (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A2 (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__I (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__I0 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A3 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A3 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__I0 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A4 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__B1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A4 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A1 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A1 (.I(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__A1 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A1 (.I(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__A1 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__A1 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A2 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__A1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__I (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__I (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__A2 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A2 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A1 (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A1 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__A2 (.I(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__A1 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__A1 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__B (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A1 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__A1 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5951__A2 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__A2 (.I(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__B2 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__A2 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__A2 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__A2 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__A2 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__B2 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__B1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__I (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A1 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__I (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__A1 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__A1 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__A1 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__A1 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__A1 (.I(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A2 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__I (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A1 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__A2 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__I (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A2 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A2 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__I (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5484__A1 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__I (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__B2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__A1 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__A2 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__I (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__A2 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__I (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__I (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A1 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A1 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__A1 (.I(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__A2 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__A2 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__A2 (.I(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A3 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__A1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__I (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__B2 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4789__I (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__B2 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__I (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__A1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__A2 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__A2 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__I (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__A2 (.I(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__A2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A2 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A2 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A2 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__A2 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__A2 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A2 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__I (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A2 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__A2 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__I (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__A3 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__B1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__A2 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__I (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__I (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__I (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__A1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__I (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__A2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__I (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A2 (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__A2 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__A2 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__A1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__A1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__B (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A2 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__I (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__A1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A2 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__A2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A1 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__A2 (.I(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5408__A1 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A1 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__A1 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__B2 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__A3 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A2 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__A3 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A1 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A1 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A1 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A1 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__I (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__I (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__I (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__B1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__A2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__I (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A2 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A2 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A2 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__A1 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A1 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__I (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__I (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__I (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__I (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A1 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__A4 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__B1 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__A1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__A2 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A2 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__I (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__B2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__I (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A1 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__A2 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A2 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__A1 (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__I (.I(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A2 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__A2 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__I (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__A1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A3 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__B1 (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__A1 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4884__I (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4867__I (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__A1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__B1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__B (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__I (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__B2 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A2 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__I (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A2 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__A3 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__A2 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__A1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__A1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__B2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A2 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__B2 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__A1 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__I (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3620__A1 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3405__A1 (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__A1 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A3 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A3 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A2 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__B1 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__B1 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__I (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__B1 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__B1 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__A1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__I (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__A3 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3405__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__A2 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__A2 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A2 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__A1 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__A1 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__A2 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3412__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__A1 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__I (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A1 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A1 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__I (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__B2 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__A1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A1 (.I(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5347__I (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__A1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__A2 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A2 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__A2 (.I(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4767__A2 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3487__A2 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3421__I (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__A1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__A2 (.I(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3408__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A2 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__A2 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4974__A1 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__A1 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__A1 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3495__A2 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__A1 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__A1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A1 (.I(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A1 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__A2 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__A2 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__A2 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__B2 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__A3 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__A2 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A2 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__I (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__A4 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__B1 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__A2 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__A1 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3788__I (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3410__A1 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A1 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__A2 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__A2 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__A1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__A2 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__A1 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3411__A2 (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__B (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__A1 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__A1 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A1 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__A2 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A3 (.I(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A2 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__I (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A1 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A2 (.I(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__A2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__A2 (.I(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__A2 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__A2 (.I(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A2 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A2 (.I(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A2 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__A2 (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__A2 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__A2 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__A2 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3626__I (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__A2 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3415__A1 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__I (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__A1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__A2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3429__I (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3415__A2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__A1 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__A2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__I (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__I0 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__I (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__I (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A2 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A1 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__A1 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__I (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__A1 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__B2 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__B2 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__I (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__B1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__A2 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__A2 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__A3 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__A1 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__A1 (.I(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__A1 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A1 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__A1 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__A1 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__A1 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__A1 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__A2 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__A1 (.I(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__I (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__B2 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__A2 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A2 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3435__A2 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3430__I (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3417__I (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5351__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__A2 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A2 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A2 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__I (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__A2 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__A1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__A1 (.I(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__A2 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A2 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__A2 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A4 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A4 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A2 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__A2 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__A1 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3428__I (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3419__I (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A2 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A2 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__A2 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__I (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__A1 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__A1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__A2 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A2 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3762__I (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3420__A2 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A1 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__A1 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__A1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__A1 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__A1 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__I (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A1 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A1 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__A1 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A2 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A2 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3688__I (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3620__A2 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__A1 (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A3 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__A1 (.I(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__A1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A2 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A2 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3708__A2 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__A2 (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3423__I (.I(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A1 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__B2 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__A1 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__A1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__A2 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A1 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__A1 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A2 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__A2 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__A2 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A2 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__A2 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3424__A2 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__A2 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__B (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__A2 (.I(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__A2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A2 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__B (.I(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__A2 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A2 (.I(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__A1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__A1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__A2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__A2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__A2 (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__A2 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__I (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A1 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__A1 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__B2 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__A1 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__I (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3426__I (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A2 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A2 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A2 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__A2 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__A2 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__B1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__A2 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A1 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__I (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__B1 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A2 (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__I (.I(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A2 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__A4 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__B2 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A2 (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__A4 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__B1 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A2 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3427__I (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__A1 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__I (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A1 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__A1 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__A2 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A2 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__A2 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__I (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__I (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__A1 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A2 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__I (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A2 (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__A2 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__A1 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__A1 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__A1 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__A2 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__A2 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__A1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__A2 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__A1 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__A2 (.I(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__A1 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A1 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__A3 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A3 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__I1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A2 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__A1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__I (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A1 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__A2 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5098__A2 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A2 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__A2 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__A2 (.I(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__A1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A1 (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__A2 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A2 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__A1 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__A1 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__A1 (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A2 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__A2 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3472__A2 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__B1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__I1 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__A2 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__A2 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A2 (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__B2 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__B1 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__A2 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__I (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__I1 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A2 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__B1 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__B1 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__A2 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__A2 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A4 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__A1 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__B1 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__A1 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A2 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__A1 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__A3 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A2 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A2 (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3431__I (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__I1 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A2 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A2 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A2 (.I(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__I (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__A2 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A2 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__A2 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3829__I (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3823__I (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3432__B2 (.I(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__A2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A2 (.I(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__B (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5172__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3433__B2 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5176__A2 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__A2 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__A1 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6785__I0 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__B2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__B2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A1 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__I (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6783__I0 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__A2 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__A2 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A2 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__A1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A1 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__A2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__A2 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__A1 (.I(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__A2 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__A2 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A3 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__A2 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__A2 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3473__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3439__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__A1 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__I (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A1 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A1 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__A2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__I (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__A1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A1 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__A1 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__A3 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__A1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__A2 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__I (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__B2 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A1 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__A1 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__A1 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A2 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__A3 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__A2 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A1 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__A2 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__A1 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__A1 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__A1 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A2 (.I(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A2 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__A2 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__A2 (.I(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4314__A2 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__I (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__A1 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3438__A2 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__A2 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__A2 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__A2 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__A2 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__A2 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__A2 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__A3 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A3 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__A2 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__A2 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3441__A2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3440__A2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__A2 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__A2 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__A3 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__A2 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__A2 (.I(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5311__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A1 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__A1 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__A2 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__A2 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__A2 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__A3 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A3 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__A3 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A1 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A2 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__A2 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__A2 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3508__A1 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3493__A1 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__I1 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A2 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__A4 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A2 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__A2 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__A2 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__A2 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A2 (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__B (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3650__I (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__A2 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3523__I (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__A2 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__A2 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__A2 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5292__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__A2 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3801__I (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3546__A2 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3445__A2 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3599__A2 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__A1 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__A1 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__B (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A4 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__B1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__A1 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__A1 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A2 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__A2 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__A2 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A3 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A2 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3799__A2 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__A2 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3448__A2 (.I(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__A1 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__A1 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__A2 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__A1 (.I(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A1 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__I (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__I (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__A1 (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3454__A2 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3449__A2 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__I1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__A2 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A2 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A2 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__A2 (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__A2 (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__A1 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A1 (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A1 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__A1 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A2 (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__I (.I(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__B2 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__A1 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A2 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__I (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A1 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__I (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3580__A1 (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3451__I (.I(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6068__A1 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__A1 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A2 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__I (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__A1 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__A1 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A2 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4291__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__A2 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__A1 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__A1 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__I (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__A2 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A2 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__A1 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6753__I1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__A1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__A1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A1 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__A2 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A1 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__B (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__A2 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3848__I (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3459__I (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3453__A2 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__A1 (.I(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__A1 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A1 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__B2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3513__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3455__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6082__A2 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__A2 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A3 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__A2 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__A2 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__A2 (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__B2 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6798__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6560__I (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__I (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__C (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__I (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__I (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__I (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6603__C (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__C (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__B (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__B (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A1 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__C (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__B (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__I (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__A2 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__A2 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__A2 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__A1 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A1 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__A1 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A3 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5406__B2 (.I(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__A1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__B2 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__A1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__A2 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__B2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__B2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3457__I (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__A1 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__A1 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__A1 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__A1 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__A1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__A2 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__A2 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A2 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A2 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A1 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__B2 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3458__I (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5424__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__A2 (.I(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A1 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A1 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A3 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A2 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A3 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__B2 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__B2 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3770__I (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3460__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A1 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A1 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__A1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__B2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__A1 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__A2 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__A2 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__A1 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__A1 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__A2 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A2 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A2 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__B2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A1 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3463__I (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__A2 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__A2 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__A1 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__B1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__A2 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__B2 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__A3 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__B2 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__B2 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3464__I (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A1 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__A1 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A1 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A1 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__A2 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__A1 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A1 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__A2 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A2 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A2 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__A2 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__I (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__B1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3466__A1 (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A1 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__A1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A1 (.I(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__A2 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__I (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A2 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3466__A2 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A1 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__A1 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__A1 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3468__A2 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3467__A2 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__A3 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__A1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__A1 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__A1 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__A1 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A1 (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3619__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3612__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3511__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3469__C (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A2 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__A2 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__A2 (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A1 (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__B2 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A2 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3492__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3491__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__A1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__A1 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A1 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5653__A1 (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__A1 (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__B (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__A2 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A2 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__A1 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__A1 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__I (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3471__A1 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__B (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A2 (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A2 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__A2 (.I(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__A1 (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__A1 (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A1 (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__B2 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A2 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A1 (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A3 (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__I (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__A2 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A1 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A1 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__B2 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__A2 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__I (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__A2 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__A2 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__A1 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3490__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__A2 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__A2 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__A1 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A1 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__A1 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__A1 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__A1 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__B2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__I (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3477__A1 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__A1 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A1 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__A1 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A2 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A1 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__A2 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__A2 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__A3 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__A2 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3477__A2 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__A2 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__A2 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A1 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__A1 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__I (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A1 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__A1 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A1 (.I(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__A2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__A1 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3479__A2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__B (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__A1 (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__A1 (.I(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5910__A1 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A1 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__A1 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A2 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A1 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A2 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__A1 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A1 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__A1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A2 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__A1 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5902__A2 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A2 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__A3 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__A1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__A1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__A2 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__A2 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3490__A2 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__A1 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__A1 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__A1 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A1 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__A2 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__B1 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__A1 (.I(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__A1 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A1 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A1 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A2 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__I (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__B2 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__B2 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__B2 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__I (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__A1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3483__A1 (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__A2 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__A2 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A2 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__A3 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A2 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__I (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3502__I (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3483__A2 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__B (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__A2 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3496__A1 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3489__A1 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__I0 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__A1 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A1 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A1 (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__I0 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__A2 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A2 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__B2 (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__A1 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4181__A2 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__I (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3621__A2 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3485__A2 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__A1 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__I (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__A2 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A2 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__A2 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5726__A1 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A1 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A3 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__A3 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__I1 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__A2 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__A1 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__A1 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__A1 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__I (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3494__A1 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3487__A1 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__A2 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5726__A2 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__A2 (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A1 (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__A1 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A2 (.I(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__A1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__A1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__A2 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__A2 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A2 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A2 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A2 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__B (.I(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__A2 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A2 (.I(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A1 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A2 (.I(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__A3 (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__A1 (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A2 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A1 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A1 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A2 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__A2 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A2 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__A2 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A2 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A2 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__A2 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__A2 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A2 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__A2 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__A1 (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__B2 (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A2 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A1 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__A1 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__A1 (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__A2 (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__A1 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__A1 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A1 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A1 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__A2 (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__I (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__A2 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__A2 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A3 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A1 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A1 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__A1 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__I1 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A1 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A1 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__A1 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A1 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A2 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__A2 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A2 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A2 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__A2 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3499__A2 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3498__A2 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__A1 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A1 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A1 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A1 (.I(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__A1 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A1 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A2 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__A1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__A1 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__A1 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__I0 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__B1 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A3 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A1 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A2 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__A2 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A2 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A3 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A3 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A2 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__A2 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__A1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__A1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__A1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A3 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__A1 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A2 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__A2 (.I(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6575__A1 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A1 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__B2 (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__B1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__A1 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A2 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__A1 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3503__I (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A2 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A2 (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__A2 (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6604__A2 (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__A2 (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__I0 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A2 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A1 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__A1 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__I1 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A2 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A2 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__A2 (.I(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__B (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6724__I1 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__A2 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__A2 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3506__A2 (.I(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6126__A1 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A1 (.I(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A1 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__A1 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A2 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__A2 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A2 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A2 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__A2 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A3 (.I(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A2 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3507__A2 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__A1 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__A1 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__A1 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__A2 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A1 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__A1 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__A1 (.I(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A1 (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__A2 (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__A3 (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__B (.I(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A2 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A1 (.I(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__I (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A2 (.I(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A2 (.I(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__A1 (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__A1 (.I(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__I0 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__A2 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A1 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A1 (.I(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5954__A1 (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__A1 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__A1 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A1 (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__I (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__A1 (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A1 (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6813__I0 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__B2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__B1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__B (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A1 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__A2 (.I(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__A2 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__A2 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A1 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__C (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A1 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__A1 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__A1 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__A2 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__B2 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__A1 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__B (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A2 (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3588__I (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3586__A2 (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3515__I (.I(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A1 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__A1 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A1 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__A1 (.I(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__B1 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3527__I (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3517__A1 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__A2 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__A2 (.I(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__A2 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__A2 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3583__I (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3517__A2 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__A2 (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__I (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__A1 (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A1 (.I(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__I (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A1 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__B (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__A1 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__A2 (.I(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__A2 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3533__A1 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3570__A2 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3519__I (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A1 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A1 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A1 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A2 (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A2 (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A2 (.I(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A2 (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A1 (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__A1 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__A1 (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__B (.I(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A2 (.I(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4247__A1 (.I(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__B2 (.I(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__A1 (.I(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A2 (.I(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__A1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A1 (.I(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__A4 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__A2 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3579__A1 (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3521__I (.I(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__A1 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__A1 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__I1 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__A1 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__A2 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A2 (.I(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__I1 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__A2 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__A1 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__B1 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__A2 (.I(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__A2 (.I(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__A2 (.I(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3522__A2 (.I(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6794__I0 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__B1 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__A1 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__B2 (.I(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__B (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__A1 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__A2 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__A1 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A1 (.I(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A2 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__B1 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A2 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__A1 (.I(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__A1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__A1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__A2 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__A2 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A2 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__A2 (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A2 (.I(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A2 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__A1 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__I (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3525__I (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__A2 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__A2 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__B (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__B (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__I (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__B (.I(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__B (.I(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__A1 (.I(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6097__B (.I(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A2 (.I(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__A1 (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__I (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__A1 (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3526__A2 (.I(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__A1 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A1 (.I(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A1 (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__A1 (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__B (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__A1 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A2 (.I(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__I (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__B1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__A1 (.I(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__B1 (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A2 (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__B2 (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__B1 (.I(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__A1 (.I(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A1 (.I(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A1 (.I(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__A2 (.I(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6639__A1 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__C (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__B (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__I (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__A3 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__A2 (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3559__I (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3531__I (.I(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A1 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A1 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__A1 (.I(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A2 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3885__I (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__I (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3532__B2 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A1 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__A1 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__I (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__A2 (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6755__I1 (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__A1 (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__A1 (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__A1 (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__I0 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A2 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A1 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__A2 (.I(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6757__I1 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__A1 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__A1 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A2 (.I(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__I1 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A1 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A1 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A1 (.I(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A2 (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__A1 (.I(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A1 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__A2 (.I(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A1 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__B (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__A2 (.I(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A1 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__A1 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3589__I (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3535__I (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A2 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A1 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__A1 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__A1 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3537__A1 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__I1 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__A2 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A2 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__A2 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__A1 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__A2 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A2 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__A2 (.I(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A1 (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__A1 (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__A3 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__B (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__A1 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3541__A1 (.I(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__A2 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__A1 (.I(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__B2 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__A2 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__A2 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__A1 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A1 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A1 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3807__I (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__I (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3545__I (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3539__I (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6774__I1 (.I(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__A2 (.I(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A2 (.I(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__A2 (.I(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__I1 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__A1 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__C (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6240__A2 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4919__A2 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__A1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__I (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3540__A2 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__A3 (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__B (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__A1 (.I(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A2 (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A3 (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__B (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3543__A2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3542__A2 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__A1 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__A1 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__B2 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__B (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__A2 (.I(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__A2 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6543__B (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__A2 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__A1 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__A2 (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__A1 (.I(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__A2 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__A2 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__A3 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__A3 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__B (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__C (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__I (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__C (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__C (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__A1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__A1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__A1 (.I(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__I (.I(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A1 (.I(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A1 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__A1 (.I(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A1 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A2 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__A1 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A1 (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__B (.I(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A2 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__A2 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__A3 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__A2 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__A4 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__A1 (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__A2 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__A2 (.I(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A2 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__I (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__A2 (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3549__I (.I(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__A2 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A2 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__A2 (.I(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__A1 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__A2 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__A2 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A2 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__B1 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3550__A2 (.I(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__A1 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6362__A1 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6361__A1 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__B (.I(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A2 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A1 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A1 (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3552__I (.I(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A1 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__A2 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__A3 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A2 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__A1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A1 (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__A1 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__A1 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__A1 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4338__A1 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A1 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__I (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__A1 (.I(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__A2 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__A2 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A2 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__I (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__A2 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3554__A2 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__A2 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A2 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__A1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__A1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__B (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6547__A2 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__A1 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__B (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3578__A1 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3573__A1 (.I(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__I (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A2 (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__A2 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__A2 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__A3 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__A1 (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A1 (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3562__I (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__A1 (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__A1 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__A1 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__A1 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__A2 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__A2 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__A2 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__A2 (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__I (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A4 (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3558__A2 (.I(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__A1 (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__A1 (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A2 (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6491__A2 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6490__A2 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A3 (.I(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__A1 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3564__A1 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__A2 (.I(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__A1 (.I(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__A1 (.I(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__A1 (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__A1 (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__A2 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__A2 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__B (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__B (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A1 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__B (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A2 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A2 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__A2 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__A1 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__A1 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__C (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__A1 (.I(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A1 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__A1 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__A1 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A1 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6448__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__B1 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__B1 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__B2 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3561__A2 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A3 (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__B (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__B (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6496__A1 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__A1 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A2 (.I(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__A2 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A1 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__A1 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__B (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A2 (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__B2 (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__A1 (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3563__A1 (.I(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__A2 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6585__A2 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__A2 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__B2 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A2 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A1 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__A1 (.I(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__B (.I(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A2 (.I(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3577__A1 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3572__A1 (.I(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__A2 (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__B (.I(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__A2 (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__A2 (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3592__A2 (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__A1 (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A2 (.I(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__B (.I(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__B (.I(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__B1 (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__B2 (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__A2 (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A2 (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__B2 (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4871__A2 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A2 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3645__A1 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3567__A2 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__A2 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__A1 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__B (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__C (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A1 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__A3 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__A2 (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A2 (.I(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A2 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A1 (.I(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A2 (.I(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__B1 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__A2 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__B (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3571__A3 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A2 (.I(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3577__A2 (.I(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3572__A2 (.I(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A3 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__A1 (.I(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6573__A2 (.I(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__A2 (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__A2 (.I(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__A1 (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3575__A2 (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3574__A2 (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__A2 (.I(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__A1 (.I(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__A2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__A1 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__A2 (.I(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6603__A2 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__A2 (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__A3 (.I(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__B (.I(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__A2 (.I(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__A3 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__B1 (.I(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__B (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6614__A2 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6615__B (.I(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__A1 (.I(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__A3 (.I(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6614__B1 (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6622__B (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__A1 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__B1 (.I(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__A2 (.I(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__A2 (.I(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__A2 (.I(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6628__A2 (.I(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6629__B (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A1 (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__A1 (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A1 (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__A2 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__A3 (.I(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__B1 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6639__A2 (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6638__A1 (.I(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__I1 (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6781__I1 (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6761__I0 (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6646__I1 (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__A1 (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__A1 (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__A1 (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6665__S (.I(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__I (.I(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6645__I (.I(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6669__A2 (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__A2 (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__S (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6646__S (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__I1 (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6783__I1 (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6763__I0 (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__I1 (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__I1 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6785__I1 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6765__I0 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__I1 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__S (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__S (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__S (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__S (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__I1 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__I1 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__I0 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__I1 (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__I (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6809__I1 (.I(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__I1 (.I(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__I0 (.I(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__I1 (.I(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__I (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A2 (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A2 (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__A2 (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3582__I (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6811__I1 (.I(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__I1 (.I(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6772__I0 (.I(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__I1 (.I(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6663__I (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6813__I1 (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6794__I1 (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6774__I0 (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6665__I1 (.I(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6666__I (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__I1 (.I(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__I1 (.I(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6718__A1 (.I(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__A1 (.I(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A1 (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A2 (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A1 (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3584__A1 (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__I0 (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__I0 (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6703__I0 (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__I0 (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6759__A1 (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6720__A1 (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__A2 (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__S (.I(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__S (.I(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__S (.I(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__S (.I(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__I0 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6724__I0 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__I0 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__I0 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A4 (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__A4 (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A2 (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3584__A2 (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__I0 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__I0 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__I0 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__I0 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__I0 (.I(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6728__I0 (.I(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6710__I0 (.I(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6684__I0 (.I(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__I0 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__I0 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__I0 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__I0 (.I(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__S (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__S (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__S (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__S (.I(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6753__I0 (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__I0 (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__I0 (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__I0 (.I(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6755__I0 (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__I0 (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__I0 (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__I0 (.I(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__I0 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6757__I0 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__I0 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__I0 (.I(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__A1 (.I(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3597__A1 (.I(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__S (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__I (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__I (.I(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6704__I (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__I (.I(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__S (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__S (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6710__S (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__S (.I(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__I (.I(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3735__A3 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__A1 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__A2 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__I (.I(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__I (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6715__I (.I(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__I (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__A1 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__B2 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__A1 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__A1 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__I (.I(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6721__I (.I(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6728__S (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__S (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6724__S (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__S (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__A4 (.I(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__B1 (.I(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4250__A2 (.I(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__B1 (.I(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__S (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__S (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__S (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6731__S (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6732__I (.I(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A1 (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__I (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__A2 (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3590__B2 (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__I (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__I (.I(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__S (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__S (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__S (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__S (.I(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__I (.I(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__I (.I(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6747__I (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6749__I (.I(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3591__B1 (.I(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__I (.I(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6754__I (.I(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__I (.I(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__I (.I(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__I (.I(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A1 (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__A1 (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__S (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6765__S (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6763__S (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6761__S (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6762__I (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6764__I (.I(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__I (.I(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__I (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6776__S (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6774__S (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6772__S (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__S (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6771__I (.I(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__I (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6775__I (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__I (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6780__I (.I(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6782__I (.I(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__S (.I(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6794__S (.I(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6792__S (.I(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__S (.I(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__I (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6799__I (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__A2 (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__A2 (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__S (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6813__S (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6811__S (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6809__S (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A2 (.I(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__A2 (.I(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3613__A2 (.I(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__A1 (.I(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3611__A1 (.I(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__A1 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__A1 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__A1 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3601__A1 (.I(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__A1 (.I(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__B (.I(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__A1 (.I(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A1 (.I(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__B2 (.I(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__I (.I(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__A1 (.I(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A2 (.I(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__A1 (.I(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3649__I (.I(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__A2 (.I(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3644__A1 (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__A2 (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__A1 (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__A2 (.I(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A3 (.I(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A1 (.I(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__A2 (.I(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__A1 (.I(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3643__A3 (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3609__A2 (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__A3 (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__A2 (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__B (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__A2 (.I(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__A2 (.I(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__A2 (.I(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3617__B (.I(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__A1 (.I(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3680__A1 (.I(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__A1 (.I(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A1 (.I(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__A1 (.I(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__A2 (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__I (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__A1 (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__B1 (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__B2 (.I(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__A1 (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__A1 (.I(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__A1 (.I(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A1 (.I(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__I (.I(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A1 (.I(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__A2 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__A2 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__A2 (.I(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__A2 (.I(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__A2 (.I(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__B2 (.I(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__A1 (.I(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__A1 (.I(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__A1 (.I(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__A2 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A2 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__A1 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__A1 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A4 (.I(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A1 (.I(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__I (.I(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__B1 (.I(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A2 (.I(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__B2 (.I(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__A1 (.I(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__A1 (.I(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__B1 (.I(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A2 (.I(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__A2 (.I(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__A2 (.I(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A3 (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__B1 (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3771__I (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__A3 (.I(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__A2 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3696__A2 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3657__A2 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__A1 (.I(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__A1 (.I(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__A2 (.I(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__I (.I(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A2 (.I(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__B2 (.I(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__A2 (.I(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__A2 (.I(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__A2 (.I(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__A2 (.I(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3714__A2 (.I(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__A2 (.I(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__A2 (.I(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3675__A2 (.I(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__A2 (.I(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__A2 (.I(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__A2 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3677__A2 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__A1 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3745__A1 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A1 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__A1 (.I(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A1 (.I(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__A2 (.I(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A2 (.I(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A2 (.I(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__I (.I(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3690__A2 (.I(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__B (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__A1 (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__A1 (.I(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3787__A1 (.I(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__A2 (.I(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__A2 (.I(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__A2 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__A1 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3705__A4 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__B1 (.I(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__A1 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__A1 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3768__A2 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__A2 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__A2 (.I(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3712__A2 (.I(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__A1 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__I (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__A1 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__A1 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A2 (.I(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A1 (.I(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__I (.I(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3723__A3 (.I(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__A1 (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3738__A1 (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A1 (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__A2 (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3731__A3 (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__I (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__A1 (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__A1 (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3735__A1 (.I(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__A2 (.I(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4226__A2 (.I(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__A2 (.I(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3735__A2 (.I(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3796__A2 (.I(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A2 (.I(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__A2 (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__A2 (.I(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__A2 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3740__A2 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3753__A2 (.I(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__A2 (.I(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__A2 (.I(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3745__A2 (.I(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__A2 (.I(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4059__A1 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__A1 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3909__A3 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__A1 (.I(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__I (.I(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__A1 (.I(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__A1 (.I(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__I (.I(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A2 (.I(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__A2 (.I(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__A1 (.I(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__I (.I(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A1 (.I(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__I (.I(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A1 (.I(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__A1 (.I(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__I1 (.I(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A2 (.I(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A2 (.I(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__A2 (.I(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__A2 (.I(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__A2 (.I(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A1 (.I(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__A1 (.I(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__A1 (.I(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__A1 (.I(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__B1 (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__A2 (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__B1 (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3763__I (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A2 (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__I (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__A2 (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3764__A2 (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__A1 (.I(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__A1 (.I(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__B (.I(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A1 (.I(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__A1 (.I(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__I (.I(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__A1 (.I(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A2 (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__A1 (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__A1 (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__I (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__A2 (.I(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__A1 (.I(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__A1 (.I(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__I (.I(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6705__I1 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A1 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__A2 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__A2 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__A1 (.I(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__A1 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__A1 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__A2 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__I (.I(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A1 (.I(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A1 (.I(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__A1 (.I(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A2 (.I(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A1 (.I(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__A2 (.I(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__I (.I(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__I0 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A2 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__A2 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__A2 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__B1 (.I(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__A1 (.I(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A2 (.I(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__A1 (.I(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A1 (.I(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A1 (.I(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__B1 (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A2 (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__I (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A2 (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A2 (.I(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A1 (.I(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A1 (.I(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__A1 (.I(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A1 (.I(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__A1 (.I(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__A1 (.I(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3787__A2 (.I(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__I (.I(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A1 (.I(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__A1 (.I(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__A1 (.I(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__A2 (.I(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A2 (.I(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3844__I (.I(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__A2 (.I(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__B1 (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__A2 (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3835__I (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3791__B1 (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3792__A2 (.I(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__A2 (.I(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__A2 (.I(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__A3 (.I(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__A1 (.I(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__A1 (.I(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A1 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__A1 (.I(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__A1 (.I(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A1 (.I(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__A2 (.I(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__A1 (.I(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A1 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3872__I (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3849__A2 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__A2 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A2 (.I(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__A2 (.I(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__A1 (.I(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__A1 (.I(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A2 (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A1 (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4114__I (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__A1 (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__A1 (.I(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A1 (.I(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__A2 (.I(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__A2 (.I(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__A2 (.I(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__A2 (.I(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3817__A2 (.I(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A2 (.I(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__A2 (.I(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4060__A1 (.I(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3821__B (.I(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__A1 (.I(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A1 (.I(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__A2 (.I(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__A1 (.I(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__A1 (.I(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A2 (.I(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__B2 (.I(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__A1 (.I(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A2 (.I(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A1 (.I(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A1 (.I(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__I (.I(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__A2 (.I(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__A2 (.I(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__A1 (.I(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__A2 (.I(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3925__A3 (.I(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__B1 (.I(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__B1 (.I(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__B1 (.I(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3912__I (.I(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3830__A2 (.I(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__A1 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__A1 (.I(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3833__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A1 (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3916__A1 (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__I (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A1 (.I(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__I (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A4 (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__B2 (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__A2 (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3919__I (.I(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__A2 (.I(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A1 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__A2 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__I (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__A2 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__A2 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__A2 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__A1 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__I (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__I (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__A1 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__A1 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__A1 (.I(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__A1 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3933__I (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__A2 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__I (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__A1 (.I(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__A2 (.I(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__I (.I(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__A2 (.I(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3960__A1 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__A1 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__A2 (.I(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__A1 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A1 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__A3 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__A3 (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__A1 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__A2 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__A1 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__A2 (.I(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__A1 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__A1 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__A1 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A1 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__I (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__I1 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A2 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A1 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__A2 (.I(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3902__A2 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__A2 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A1 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__A1 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__A1 (.I(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3895__A1 (.I(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__I1 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A2 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__B1 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__A2 (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__I (.I(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__I1 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__B1 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__A2 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__B1 (.I(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A2 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__B2 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__I (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__B2 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__A2 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__A2 (.I(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__B1 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__A1 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3935__I (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3878__A1 (.I(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__A2 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__A1 (.I(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__B2 (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__B2 (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__A1 (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__A1 (.I(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3951__A3 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__B1 (.I(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A2 (.I(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A1 (.I(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__A2 (.I(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A1 (.I(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__A1 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__B2 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__I (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__B2 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__A1 (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__A1 (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__A1 (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3962__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3890__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__A2 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__A1 (.I(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__A1 (.I(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__A2 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__A2 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A2 (.I(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__A2 (.I(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__B (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A2 (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__A2 (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__A1 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4055__A1 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__B1 (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__A2 (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__I (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__A2 (.I(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__I0 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__A2 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__A1 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3916__A2 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3931__A2 (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3929__A1 (.I(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3925__A2 (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__A1 (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__A1 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__A2 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__B2 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__A1 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__A1 (.I(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__A2 (.I(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__A1 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__A1 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__A2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__A2 (.I(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__A2 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__I (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A1 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3934__A1 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__A2 (.I(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4534__A1 (.I(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__I (.I(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__A2 (.I(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__A1 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__A1 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__A3 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6765__I1 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__A2 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__A2 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__A2 (.I(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4008__A1 (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__A1 (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__A2 (.I(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A1 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__I (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__A1 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__A1 (.I(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6703__I1 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A1 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__A1 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__A2 (.I(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__A1 (.I(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A1 (.I(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__A2 (.I(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__A3 (.I(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__A1 (.I(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A1 (.I(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__A1 (.I(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A2 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__A2 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A1 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__A2 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__A1 (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__A1 (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__A2 (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__A2 (.I(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A2 (.I(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4086__I (.I(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__B1 (.I(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__A1 (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__A1 (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__A2 (.I(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__A2 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__A2 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__A3 (.I(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__A2 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A2 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__A2 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__A1 (.I(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__A1 (.I(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__A1 (.I(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__I (.I(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__A2 (.I(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__A2 (.I(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__A2 (.I(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3973__A1 (.I(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__A1 (.I(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3964__A2 (.I(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__A2 (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__A2 (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3965__A2 (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A1 (.I(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A1 (.I(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__A2 (.I(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A2 (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A2 (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__A3 (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A3 (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__A2 (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A2 (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A1 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__A1 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__A2 (.I(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3989__A2 (.I(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A3 (.I(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A2 (.I(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__A2 (.I(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__A1 (.I(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__A1 (.I(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A1 (.I(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A2 (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4048__A2 (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A3 (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__A2 (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__A1 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__A1 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__A3 (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4005__A1 (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4036__A2 (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__A2 (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A1 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__A1 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6763__I1 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A2 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A4 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__A2 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__A2 (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__A2 (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A1 (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__A2 (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__A2 (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__I0 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4657__A2 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A2 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A2 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A1 (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__A1 (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A2 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__A2 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A1 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A1 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A2 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__I (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A1 (.I(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A1 (.I(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__I (.I(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__A1 (.I(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__A1 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A3 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__A3 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A1 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4031__A1 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A2 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__A2 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6538__A1 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__A2 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4043__A2 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4040__A3 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A1 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A1 (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A1 (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A1 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__A1 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__A2 (.I(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__A1 (.I(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__A1 (.I(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4047__A2 (.I(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6596__A2 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__B2 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6615__A1 (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__B2 (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__A1 (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6615__A2 (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__B3 (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__A2 (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__A3 (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A2 (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__A2 (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__A1 (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A1 (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__A1 (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__B (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__A1 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__A2 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A1 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A1 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__A1 (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__A1 (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__A1 (.I(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6728__I1 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__A2 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A2 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__A2 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__A1 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__A1 (.I(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__I (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__A1 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__A2 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A1 (.I(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A2 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A3 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__B1 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4085__I (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__I (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__A2 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__A2 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A2 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__I1 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A3 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__A2 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A3 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6710__I1 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A4 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__B1 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4088__A4 (.I(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__A1 (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__A1 (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__A2 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__I (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__A1 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A1 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A2 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__A2 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__A1 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A1 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__A2 (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A1 (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__A1 (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__A1 (.I(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6772__I1 (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A2 (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A1 (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4105__A1 (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__A2 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A1 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A1 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__I (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__A1 (.I(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A1 (.I(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__B1 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__A2 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A4 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4112__I (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A2 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A1 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__B2 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A1 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__A1 (.I(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A1 (.I(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4116__A2 (.I(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__A2 (.I(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4119__A2 (.I(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A2 (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__A2 (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A3 (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__A2 (.I(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__A2 (.I(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4127__A2 (.I(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A3 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__A2 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__A2 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__A2 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__I (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__I (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__A2 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__A1 (.I(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__A1 (.I(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A1 (.I(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__I (.I(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__A1 (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__A1 (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__B (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A1 (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A1 (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A1 (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__I (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A2 (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A2 (.I(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A1 (.I(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__I (.I(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__A1 (.I(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__I (.I(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__I (.I(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__A2 (.I(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__A2 (.I(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__A2 (.I(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__A1 (.I(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__B2 (.I(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A1 (.I(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__A2 (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__I (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A2 (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__I (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__A2 (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__A2 (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__A2 (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A2 (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A2 (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__I (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__A2 (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A1 (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A2 (.I(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__B1 (.I(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__A2 (.I(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__B1 (.I(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A3 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__A2 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A2 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__A1 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__A1 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A1 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__A1 (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A3 (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__I (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A1 (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__A1 (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__A1 (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A1 (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__A1 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__A2 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A2 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A1 (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A2 (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__A2 (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4169__A2 (.I(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__A1 (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__A1 (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4382__A2 (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__I (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__I (.I(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A2 (.I(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__A1 (.I(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4175__A1 (.I(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A1 (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A1 (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__A1 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A1 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__A1 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4187__A1 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A1 (.I(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__B2 (.I(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__A1 (.I(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A1 (.I(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__A2 (.I(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__I (.I(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__A2 (.I(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__A2 (.I(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A2 (.I(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__A2 (.I(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__A2 (.I(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__A2 (.I(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__B2 (.I(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__A1 (.I(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__B2 (.I(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__I (.I(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__B1 (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A1 (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__B1 (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__I (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__I (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A1 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A1 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__A3 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A1 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__A2 (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__A2 (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__I (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__I (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__B2 (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A4 (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__I (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__A2 (.I(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A2 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4325__I (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4243__A1 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4223__I (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A2 (.I(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__I (.I(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__B1 (.I(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4226__A1 (.I(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__A2 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5437__A2 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__B2 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__B1 (.I(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A1 (.I(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4236__A1 (.I(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A2 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__A2 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4449__A3 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__A2 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__I (.I(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A1 (.I(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A1 (.I(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__I (.I(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A1 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__B2 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__I (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A1 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A2 (.I(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4236__A2 (.I(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A1 (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__I (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__I (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4240__A1 (.I(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(execute));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(input_val[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(input_val[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(input_val[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(input_val[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(input_val[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(input_val[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(input_val[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(input_val[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(reset));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(sel_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(sel_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(sel_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(sel_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(sel_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6880__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6871__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6870__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6863__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6862__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6855__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6854__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6853__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6846__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6842__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6835__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6825__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6819__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6818__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6641__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6648__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6651__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6686__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6658__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6690__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6693__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6880__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6879__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6871__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6870__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6869__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6863__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6862__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6855__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6854__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6853__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6851__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6846__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6845__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6842__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6841__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6839__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6835__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6825__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6822__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6819__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6818__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__RN (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6779__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__A2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__A2 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6778__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3400__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3401__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output17_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output19_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output23_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1223 ();
endmodule

